/*
 
 Conway's Game of Life modeled in SVerilog
 
 */

module datapath ( grid, grid_evolve );

   output logic [1023:0] 	grid_evolve;
   input logic [1023:0] 	grid;
   


evolve3 e0 (grid_evolve[0], grid[1], grid[32], grid[33], grid[0]);
evolve5 e1 (grid_evolve[1], grid[0], grid[2], grid[32], grid[33], grid[34], grid[1]);
evolve5 e2 (grid_evolve[2], grid[1], grid[3], grid[33], grid[34], grid[35], grid[2]);
evolve5 e3 (grid_evolve[3], grid[2], grid[4], grid[34], grid[35], grid[36], grid[3]);
evolve5 e4 (grid_evolve[4], grid[3], grid[5], grid[35], grid[36], grid[37], grid[4]);
evolve5 e5 (grid_evolve[5], grid[4], grid[6], grid[36], grid[37], grid[38], grid[5]);
evolve5 e6 (grid_evolve[6], grid[5], grid[7], grid[37], grid[38], grid[39], grid[6]);
evolve5 e7 (grid_evolve[7], grid[6], grid[8], grid[38], grid[39], grid[40], grid[7]);
evolve5 e8 (grid_evolve[8], grid[7], grid[9], grid[39], grid[40], grid[41], grid[8]);
evolve5 e9 (grid_evolve[9], grid[8], grid[10], grid[40], grid[41], grid[42], grid[9]);
evolve5 e10 (grid_evolve[10], grid[9], grid[11], grid[41], grid[42], grid[43], grid[10]);
evolve5 e11 (grid_evolve[11], grid[10], grid[12], grid[42], grid[43], grid[44], grid[11]);
evolve5 e12 (grid_evolve[12], grid[11], grid[13], grid[43], grid[44], grid[45], grid[12]);
evolve5 e13 (grid_evolve[13], grid[12], grid[14], grid[44], grid[45], grid[46], grid[13]);
evolve5 e14 (grid_evolve[14], grid[13], grid[15], grid[45], grid[46], grid[47], grid[14]);
evolve5 e15 (grid_evolve[15], grid[14], grid[16], grid[46], grid[47], grid[48], grid[15]);
evolve5 e16 (grid_evolve[16], grid[15], grid[17], grid[47], grid[48], grid[49], grid[16]);
evolve5 e17 (grid_evolve[17], grid[16], grid[18], grid[48], grid[49], grid[50], grid[17]);
evolve5 e18 (grid_evolve[18], grid[17], grid[19], grid[49], grid[50], grid[51], grid[18]);
evolve5 e19 (grid_evolve[19], grid[18], grid[20], grid[50], grid[51], grid[52], grid[19]);
evolve5 e20 (grid_evolve[20], grid[19], grid[21], grid[51], grid[52], grid[53], grid[20]);
evolve5 e21 (grid_evolve[21], grid[20], grid[22], grid[52], grid[53], grid[54], grid[21]);
evolve5 e22 (grid_evolve[22], grid[21], grid[23], grid[53], grid[54], grid[55], grid[22]);
evolve5 e23 (grid_evolve[23], grid[22], grid[24], grid[54], grid[55], grid[56], grid[23]);
evolve5 e24 (grid_evolve[24], grid[23], grid[25], grid[55], grid[56], grid[57], grid[24]);
evolve5 e25 (grid_evolve[25], grid[24], grid[26], grid[56], grid[57], grid[58], grid[25]);
evolve5 e26 (grid_evolve[26], grid[25], grid[27], grid[57], grid[58], grid[59], grid[26]);
evolve5 e27 (grid_evolve[27], grid[26], grid[28], grid[58], grid[59], grid[60], grid[27]);
evolve5 e28 (grid_evolve[28], grid[27], grid[29], grid[59], grid[60], grid[61], grid[28]);
evolve5 e29 (grid_evolve[29], grid[28], grid[30], grid[60], grid[61], grid[62], grid[29]);
evolve5 e30 (grid_evolve[30], grid[29], grid[31], grid[61], grid[62], grid[63], grid[30]);
evolve3 e31 (grid_evolve[31], grid[30], grid[62], grid[63], grid[31]);

evolve5 e32 (grid_evolve[32], grid[0], grid[1], grid[33], grid[64], grid[65], grid[32]);
evolve8 e33 (grid_evolve[33], grid[0], grid[1], grid[2], grid[32], grid[34], grid[64], grid[65], grid[66], grid[33]);
evolve8 e34 (grid_evolve[34], grid[1], grid[2], grid[3], grid[33], grid[35], grid[65], grid[66], grid[67], grid[34]);
evolve8 e35 (grid_evolve[35], grid[2], grid[3], grid[4], grid[34], grid[36], grid[66], grid[67], grid[68], grid[35]);
evolve8 e36 (grid_evolve[36], grid[3], grid[4], grid[5], grid[35], grid[37], grid[67], grid[68], grid[69], grid[36]);
evolve8 e37 (grid_evolve[37], grid[4], grid[5], grid[6], grid[36], grid[38], grid[68], grid[69], grid[70], grid[37]);
evolve8 e38 (grid_evolve[38], grid[5], grid[6], grid[7], grid[37], grid[39], grid[69], grid[70], grid[71], grid[38]);
evolve8 e39 (grid_evolve[39], grid[6], grid[7], grid[8], grid[38], grid[40], grid[70], grid[71], grid[72], grid[39]);
evolve8 e40 (grid_evolve[40], grid[7], grid[8], grid[9], grid[39], grid[41], grid[71], grid[72], grid[73], grid[40]);
evolve8 e41 (grid_evolve[41], grid[8], grid[9], grid[10], grid[40], grid[42], grid[72], grid[73], grid[74], grid[41]);
evolve8 e42 (grid_evolve[42], grid[9], grid[10], grid[11], grid[41], grid[43], grid[73], grid[74], grid[75], grid[42]);
evolve8 e43 (grid_evolve[43], grid[10], grid[11], grid[12], grid[42], grid[44], grid[74], grid[75], grid[76], grid[43]);
evolve8 e44 (grid_evolve[44], grid[11], grid[12], grid[13], grid[43], grid[45], grid[75], grid[76], grid[77], grid[44]);
evolve8 e45 (grid_evolve[45], grid[12], grid[13], grid[14], grid[44], grid[46], grid[76], grid[77], grid[78], grid[45]);
evolve8 e46 (grid_evolve[46], grid[13], grid[14], grid[15], grid[45], grid[47], grid[77], grid[78], grid[79], grid[46]);
evolve8 e47 (grid_evolve[47], grid[14], grid[15], grid[16], grid[46], grid[48], grid[78], grid[79], grid[80], grid[47]);
evolve8 e48 (grid_evolve[48], grid[15], grid[16], grid[17], grid[47], grid[49], grid[79], grid[80], grid[81], grid[48]);
evolve8 e49 (grid_evolve[49], grid[16], grid[17], grid[18], grid[48], grid[50], grid[80], grid[81], grid[82], grid[49]);
evolve8 e50 (grid_evolve[50], grid[17], grid[18], grid[19], grid[49], grid[51], grid[81], grid[82], grid[83], grid[50]);
evolve8 e51 (grid_evolve[51], grid[18], grid[19], grid[20], grid[50], grid[52], grid[82], grid[83], grid[84], grid[51]);
evolve8 e52 (grid_evolve[52], grid[19], grid[20], grid[21], grid[51], grid[53], grid[83], grid[84], grid[85], grid[52]);
evolve8 e53 (grid_evolve[53], grid[20], grid[21], grid[22], grid[52], grid[54], grid[84], grid[85], grid[86], grid[53]);
evolve8 e54 (grid_evolve[54], grid[21], grid[22], grid[23], grid[53], grid[55], grid[85], grid[86], grid[87], grid[54]);
evolve8 e55 (grid_evolve[55], grid[22], grid[23], grid[24], grid[54], grid[56], grid[86], grid[87], grid[88], grid[55]);
evolve8 e56 (grid_evolve[56], grid[23], grid[24], grid[25], grid[55], grid[57], grid[87], grid[88], grid[89], grid[56]);
evolve8 e57 (grid_evolve[57], grid[24], grid[25], grid[26], grid[56], grid[58], grid[88], grid[89], grid[90], grid[57]);
evolve8 e58 (grid_evolve[58], grid[25], grid[26], grid[27], grid[57], grid[59], grid[89], grid[90], grid[91], grid[58]);
evolve8 e59 (grid_evolve[59], grid[26], grid[27], grid[28], grid[58], grid[60], grid[90], grid[91], grid[92], grid[59]);
evolve8 e60 (grid_evolve[60], grid[27], grid[28], grid[29], grid[59], grid[61], grid[91], grid[92], grid[93], grid[60]);
evolve8 e61 (grid_evolve[61], grid[28], grid[29], grid[30], grid[60], grid[62], grid[92], grid[93], grid[94], grid[61]);
evolve8 e62 (grid_evolve[62], grid[29], grid[30], grid[31], grid[61], grid[63], grid[93], grid[94], grid[95], grid[62]);
evolve5 e63 (grid_evolve[63], grid[30], grid[31], grid[62], grid[94], grid[95], grid[63]);

evolve5 e64 (grid_evolve[64], grid[32], grid[33], grid[65], grid[96], grid[97], grid[64]);
evolve8 e65 (grid_evolve[65], grid[32], grid[33], grid[34], grid[64], grid[66], grid[96], grid[97], grid[98], grid[65]);
evolve8 e66 (grid_evolve[66], grid[33], grid[34], grid[35], grid[65], grid[67], grid[97], grid[98], grid[99], grid[66]);
evolve8 e67 (grid_evolve[67], grid[34], grid[35], grid[36], grid[66], grid[68], grid[98], grid[99], grid[100], grid[67]);
evolve8 e68 (grid_evolve[68], grid[35], grid[36], grid[37], grid[67], grid[69], grid[99], grid[100], grid[101], grid[68]);
evolve8 e69 (grid_evolve[69], grid[36], grid[37], grid[38], grid[68], grid[70], grid[100], grid[101], grid[102], grid[69]);
evolve8 e70 (grid_evolve[70], grid[37], grid[38], grid[39], grid[69], grid[71], grid[101], grid[102], grid[103], grid[70]);
evolve8 e71 (grid_evolve[71], grid[38], grid[39], grid[40], grid[70], grid[72], grid[102], grid[103], grid[104], grid[71]);
evolve8 e72 (grid_evolve[72], grid[39], grid[40], grid[41], grid[71], grid[73], grid[103], grid[104], grid[105], grid[72]);
evolve8 e73 (grid_evolve[73], grid[40], grid[41], grid[42], grid[72], grid[74], grid[104], grid[105], grid[106], grid[73]);
evolve8 e74 (grid_evolve[74], grid[41], grid[42], grid[43], grid[73], grid[75], grid[105], grid[106], grid[107], grid[74]);
evolve8 e75 (grid_evolve[75], grid[42], grid[43], grid[44], grid[74], grid[76], grid[106], grid[107], grid[108], grid[75]);
evolve8 e76 (grid_evolve[76], grid[43], grid[44], grid[45], grid[75], grid[77], grid[107], grid[108], grid[109], grid[76]);
evolve8 e77 (grid_evolve[77], grid[44], grid[45], grid[46], grid[76], grid[78], grid[108], grid[109], grid[110], grid[77]);
evolve8 e78 (grid_evolve[78], grid[45], grid[46], grid[47], grid[77], grid[79], grid[109], grid[110], grid[111], grid[78]);
evolve8 e79 (grid_evolve[79], grid[46], grid[47], grid[48], grid[78], grid[80], grid[110], grid[111], grid[112], grid[79]);
evolve8 e80 (grid_evolve[80], grid[47], grid[48], grid[49], grid[79], grid[81], grid[111], grid[112], grid[113], grid[80]);
evolve8 e81 (grid_evolve[81], grid[48], grid[49], grid[50], grid[80], grid[82], grid[112], grid[113], grid[114], grid[81]);
evolve8 e82 (grid_evolve[82], grid[49], grid[50], grid[51], grid[81], grid[83], grid[113], grid[114], grid[115], grid[82]);
evolve8 e83 (grid_evolve[83], grid[50], grid[51], grid[52], grid[82], grid[84], grid[114], grid[115], grid[116], grid[83]);
evolve8 e84 (grid_evolve[84], grid[51], grid[52], grid[53], grid[83], grid[85], grid[115], grid[116], grid[117], grid[84]);
evolve8 e85 (grid_evolve[85], grid[52], grid[53], grid[54], grid[84], grid[86], grid[116], grid[117], grid[118], grid[85]);
evolve8 e86 (grid_evolve[86], grid[53], grid[54], grid[55], grid[85], grid[87], grid[117], grid[118], grid[119], grid[86]);
evolve8 e87 (grid_evolve[87], grid[54], grid[55], grid[56], grid[86], grid[88], grid[118], grid[119], grid[120], grid[87]);
evolve8 e88 (grid_evolve[88], grid[55], grid[56], grid[57], grid[87], grid[89], grid[119], grid[120], grid[121], grid[88]);
evolve8 e89 (grid_evolve[89], grid[56], grid[57], grid[58], grid[88], grid[90], grid[120], grid[121], grid[122], grid[89]);
evolve8 e90 (grid_evolve[90], grid[57], grid[58], grid[59], grid[89], grid[91], grid[121], grid[122], grid[123], grid[90]);
evolve8 e91 (grid_evolve[91], grid[58], grid[59], grid[60], grid[90], grid[92], grid[122], grid[123], grid[124], grid[91]);
evolve8 e92 (grid_evolve[92], grid[59], grid[60], grid[61], grid[91], grid[93], grid[123], grid[124], grid[125], grid[92]);
evolve8 e93 (grid_evolve[93], grid[60], grid[61], grid[62], grid[92], grid[94], grid[124], grid[125], grid[126], grid[93]);
evolve8 e94 (grid_evolve[94], grid[61], grid[62], grid[63], grid[93], grid[95], grid[125], grid[126], grid[127], grid[94]);
evolve5 e95 (grid_evolve[95], grid[62], grid[63], grid[94], grid[126], grid[127], grid[95]);

evolve5 e96 (grid_evolve[96], grid[64], grid[65], grid[97], grid[128], grid[129], grid[96]);
evolve8 e97 (grid_evolve[97], grid[64], grid[65], grid[66], grid[96], grid[98], grid[128], grid[129], grid[130], grid[97]);
evolve8 e98 (grid_evolve[98], grid[65], grid[66], grid[67], grid[97], grid[99], grid[129], grid[130], grid[131], grid[98]);
evolve8 e99 (grid_evolve[99], grid[66], grid[67], grid[68], grid[98], grid[100], grid[130], grid[131], grid[132], grid[99]);
evolve8 e100 (grid_evolve[100], grid[67], grid[68], grid[69], grid[99], grid[101], grid[131], grid[132], grid[133], grid[100]);
evolve8 e101 (grid_evolve[101], grid[68], grid[69], grid[70], grid[100], grid[102], grid[132], grid[133], grid[134], grid[101]);
evolve8 e102 (grid_evolve[102], grid[69], grid[70], grid[71], grid[101], grid[103], grid[133], grid[134], grid[135], grid[102]);
evolve8 e103 (grid_evolve[103], grid[70], grid[71], grid[72], grid[102], grid[104], grid[134], grid[135], grid[136], grid[103]);
evolve8 e104 (grid_evolve[104], grid[71], grid[72], grid[73], grid[103], grid[105], grid[135], grid[136], grid[137], grid[104]);
evolve8 e105 (grid_evolve[105], grid[72], grid[73], grid[74], grid[104], grid[106], grid[136], grid[137], grid[138], grid[105]);
evolve8 e106 (grid_evolve[106], grid[73], grid[74], grid[75], grid[105], grid[107], grid[137], grid[138], grid[139], grid[106]);
evolve8 e107 (grid_evolve[107], grid[74], grid[75], grid[76], grid[106], grid[108], grid[138], grid[139], grid[140], grid[107]);
evolve8 e108 (grid_evolve[108], grid[75], grid[76], grid[77], grid[107], grid[109], grid[139], grid[140], grid[141], grid[108]);
evolve8 e109 (grid_evolve[109], grid[76], grid[77], grid[78], grid[108], grid[110], grid[140], grid[141], grid[142], grid[109]);
evolve8 e110 (grid_evolve[110], grid[77], grid[78], grid[79], grid[109], grid[111], grid[141], grid[142], grid[143], grid[110]);
evolve8 e111 (grid_evolve[111], grid[78], grid[79], grid[80], grid[110], grid[112], grid[142], grid[143], grid[144], grid[111]);
evolve8 e112 (grid_evolve[112], grid[79], grid[80], grid[81], grid[111], grid[113], grid[143], grid[144], grid[145], grid[112]);
evolve8 e113 (grid_evolve[113], grid[80], grid[81], grid[82], grid[112], grid[114], grid[144], grid[145], grid[146], grid[113]);
evolve8 e114 (grid_evolve[114], grid[81], grid[82], grid[83], grid[113], grid[115], grid[145], grid[146], grid[147], grid[114]);
evolve8 e115 (grid_evolve[115], grid[82], grid[83], grid[84], grid[114], grid[116], grid[146], grid[147], grid[148], grid[115]);
evolve8 e116 (grid_evolve[116], grid[83], grid[84], grid[85], grid[115], grid[117], grid[147], grid[148], grid[149], grid[116]);
evolve8 e117 (grid_evolve[117], grid[84], grid[85], grid[86], grid[116], grid[118], grid[148], grid[149], grid[150], grid[117]);
evolve8 e118 (grid_evolve[118], grid[85], grid[86], grid[87], grid[117], grid[119], grid[149], grid[150], grid[151], grid[118]);
evolve8 e119 (grid_evolve[119], grid[86], grid[87], grid[88], grid[118], grid[120], grid[150], grid[151], grid[152], grid[119]);
evolve8 e120 (grid_evolve[120], grid[87], grid[88], grid[89], grid[119], grid[121], grid[151], grid[152], grid[153], grid[120]);
evolve8 e121 (grid_evolve[121], grid[88], grid[89], grid[90], grid[120], grid[122], grid[152], grid[153], grid[154], grid[121]);
evolve8 e122 (grid_evolve[122], grid[89], grid[90], grid[91], grid[121], grid[123], grid[153], grid[154], grid[155], grid[122]);
evolve8 e123 (grid_evolve[123], grid[90], grid[91], grid[92], grid[122], grid[124], grid[154], grid[155], grid[156], grid[123]);
evolve8 e124 (grid_evolve[124], grid[91], grid[92], grid[93], grid[123], grid[125], grid[155], grid[156], grid[157], grid[124]);
evolve8 e125 (grid_evolve[125], grid[92], grid[93], grid[94], grid[124], grid[126], grid[156], grid[157], grid[158], grid[125]);
evolve8 e126 (grid_evolve[126], grid[93], grid[94], grid[95], grid[125], grid[127], grid[157], grid[158], grid[159], grid[126]);
evolve5 e127 (grid_evolve[127], grid[94], grid[95], grid[126], grid[158], grid[159], grid[127]);

evolve5 e128 (grid_evolve[128], grid[96], grid[97], grid[129], grid[160], grid[161], grid[128]);
evolve8 e129 (grid_evolve[129], grid[96], grid[97], grid[98], grid[128], grid[130], grid[160], grid[161], grid[162], grid[129]);
evolve8 e130 (grid_evolve[130], grid[97], grid[98], grid[99], grid[129], grid[131], grid[161], grid[162], grid[163], grid[130]);
evolve8 e131 (grid_evolve[131], grid[98], grid[99], grid[100], grid[130], grid[132], grid[162], grid[163], grid[164], grid[131]);
evolve8 e132 (grid_evolve[132], grid[99], grid[100], grid[101], grid[131], grid[133], grid[163], grid[164], grid[165], grid[132]);
evolve8 e133 (grid_evolve[133], grid[100], grid[101], grid[102], grid[132], grid[134], grid[164], grid[165], grid[166], grid[133]);
evolve8 e134 (grid_evolve[134], grid[101], grid[102], grid[103], grid[133], grid[135], grid[165], grid[166], grid[167], grid[134]);
evolve8 e135 (grid_evolve[135], grid[102], grid[103], grid[104], grid[134], grid[136], grid[166], grid[167], grid[168], grid[135]);
evolve8 e136 (grid_evolve[136], grid[103], grid[104], grid[105], grid[135], grid[137], grid[167], grid[168], grid[169], grid[136]);
evolve8 e137 (grid_evolve[137], grid[104], grid[105], grid[106], grid[136], grid[138], grid[168], grid[169], grid[170], grid[137]);
evolve8 e138 (grid_evolve[138], grid[105], grid[106], grid[107], grid[137], grid[139], grid[169], grid[170], grid[171], grid[138]);
evolve8 e139 (grid_evolve[139], grid[106], grid[107], grid[108], grid[138], grid[140], grid[170], grid[171], grid[172], grid[139]);
evolve8 e140 (grid_evolve[140], grid[107], grid[108], grid[109], grid[139], grid[141], grid[171], grid[172], grid[173], grid[140]);
evolve8 e141 (grid_evolve[141], grid[108], grid[109], grid[110], grid[140], grid[142], grid[172], grid[173], grid[174], grid[141]);
evolve8 e142 (grid_evolve[142], grid[109], grid[110], grid[111], grid[141], grid[143], grid[173], grid[174], grid[175], grid[142]);
evolve8 e143 (grid_evolve[143], grid[110], grid[111], grid[112], grid[142], grid[144], grid[174], grid[175], grid[176], grid[143]);
evolve8 e144 (grid_evolve[144], grid[111], grid[112], grid[113], grid[143], grid[145], grid[175], grid[176], grid[177], grid[144]);
evolve8 e145 (grid_evolve[145], grid[112], grid[113], grid[114], grid[144], grid[146], grid[176], grid[177], grid[178], grid[145]);
evolve8 e146 (grid_evolve[146], grid[113], grid[114], grid[115], grid[145], grid[147], grid[177], grid[178], grid[179], grid[146]);
evolve8 e147 (grid_evolve[147], grid[114], grid[115], grid[116], grid[146], grid[148], grid[178], grid[179], grid[180], grid[147]);
evolve8 e148 (grid_evolve[148], grid[115], grid[116], grid[117], grid[147], grid[149], grid[179], grid[180], grid[181], grid[148]);
evolve8 e149 (grid_evolve[149], grid[116], grid[117], grid[118], grid[148], grid[150], grid[180], grid[181], grid[182], grid[149]);
evolve8 e150 (grid_evolve[150], grid[117], grid[118], grid[119], grid[149], grid[151], grid[181], grid[182], grid[183], grid[150]);
evolve8 e151 (grid_evolve[151], grid[118], grid[119], grid[120], grid[150], grid[152], grid[182], grid[183], grid[184], grid[151]);
evolve8 e152 (grid_evolve[152], grid[119], grid[120], grid[121], grid[151], grid[153], grid[183], grid[184], grid[185], grid[152]);
evolve8 e153 (grid_evolve[153], grid[120], grid[121], grid[122], grid[152], grid[154], grid[184], grid[185], grid[186], grid[153]);
evolve8 e154 (grid_evolve[154], grid[121], grid[122], grid[123], grid[153], grid[155], grid[185], grid[186], grid[187], grid[154]);
evolve8 e155 (grid_evolve[155], grid[122], grid[123], grid[124], grid[154], grid[156], grid[186], grid[187], grid[188], grid[155]);
evolve8 e156 (grid_evolve[156], grid[123], grid[124], grid[125], grid[155], grid[157], grid[187], grid[188], grid[189], grid[156]);
evolve8 e157 (grid_evolve[157], grid[124], grid[125], grid[126], grid[156], grid[158], grid[188], grid[189], grid[190], grid[157]);
evolve8 e158 (grid_evolve[158], grid[125], grid[126], grid[127], grid[157], grid[159], grid[189], grid[190], grid[191], grid[158]);
evolve5 e159 (grid_evolve[159], grid[126], grid[127], grid[158], grid[190], grid[191], grid[159]);

evolve5 e160 (grid_evolve[160], grid[128], grid[129], grid[161], grid[192], grid[193], grid[160]);
evolve8 e161 (grid_evolve[161], grid[128], grid[129], grid[130], grid[160], grid[162], grid[192], grid[193], grid[194], grid[161]);
evolve8 e162 (grid_evolve[162], grid[129], grid[130], grid[131], grid[161], grid[163], grid[193], grid[194], grid[195], grid[162]);
evolve8 e163 (grid_evolve[163], grid[130], grid[131], grid[132], grid[162], grid[164], grid[194], grid[195], grid[196], grid[163]);
evolve8 e164 (grid_evolve[164], grid[131], grid[132], grid[133], grid[163], grid[165], grid[195], grid[196], grid[197], grid[164]);
evolve8 e165 (grid_evolve[165], grid[132], grid[133], grid[134], grid[164], grid[166], grid[196], grid[197], grid[198], grid[165]);
evolve8 e166 (grid_evolve[166], grid[133], grid[134], grid[135], grid[165], grid[167], grid[197], grid[198], grid[199], grid[166]);
evolve8 e167 (grid_evolve[167], grid[134], grid[135], grid[136], grid[166], grid[168], grid[198], grid[199], grid[200], grid[167]);
evolve8 e168 (grid_evolve[168], grid[135], grid[136], grid[137], grid[167], grid[169], grid[199], grid[200], grid[201], grid[168]);
evolve8 e169 (grid_evolve[169], grid[136], grid[137], grid[138], grid[168], grid[170], grid[200], grid[201], grid[202], grid[169]);
evolve8 e170 (grid_evolve[170], grid[137], grid[138], grid[139], grid[169], grid[171], grid[201], grid[202], grid[203], grid[170]);
evolve8 e171 (grid_evolve[171], grid[138], grid[139], grid[140], grid[170], grid[172], grid[202], grid[203], grid[204], grid[171]);
evolve8 e172 (grid_evolve[172], grid[139], grid[140], grid[141], grid[171], grid[173], grid[203], grid[204], grid[205], grid[172]);
evolve8 e173 (grid_evolve[173], grid[140], grid[141], grid[142], grid[172], grid[174], grid[204], grid[205], grid[206], grid[173]);
evolve8 e174 (grid_evolve[174], grid[141], grid[142], grid[143], grid[173], grid[175], grid[205], grid[206], grid[207], grid[174]);
evolve8 e175 (grid_evolve[175], grid[142], grid[143], grid[144], grid[174], grid[176], grid[206], grid[207], grid[208], grid[175]);
evolve8 e176 (grid_evolve[176], grid[143], grid[144], grid[145], grid[175], grid[177], grid[207], grid[208], grid[209], grid[176]);
evolve8 e177 (grid_evolve[177], grid[144], grid[145], grid[146], grid[176], grid[178], grid[208], grid[209], grid[210], grid[177]);
evolve8 e178 (grid_evolve[178], grid[145], grid[146], grid[147], grid[177], grid[179], grid[209], grid[210], grid[211], grid[178]);
evolve8 e179 (grid_evolve[179], grid[146], grid[147], grid[148], grid[178], grid[180], grid[210], grid[211], grid[212], grid[179]);
evolve8 e180 (grid_evolve[180], grid[147], grid[148], grid[149], grid[179], grid[181], grid[211], grid[212], grid[213], grid[180]);
evolve8 e181 (grid_evolve[181], grid[148], grid[149], grid[150], grid[180], grid[182], grid[212], grid[213], grid[214], grid[181]);
evolve8 e182 (grid_evolve[182], grid[149], grid[150], grid[151], grid[181], grid[183], grid[213], grid[214], grid[215], grid[182]);
evolve8 e183 (grid_evolve[183], grid[150], grid[151], grid[152], grid[182], grid[184], grid[214], grid[215], grid[216], grid[183]);
evolve8 e184 (grid_evolve[184], grid[151], grid[152], grid[153], grid[183], grid[185], grid[215], grid[216], grid[217], grid[184]);
evolve8 e185 (grid_evolve[185], grid[152], grid[153], grid[154], grid[184], grid[186], grid[216], grid[217], grid[218], grid[185]);
evolve8 e186 (grid_evolve[186], grid[153], grid[154], grid[155], grid[185], grid[187], grid[217], grid[218], grid[219], grid[186]);
evolve8 e187 (grid_evolve[187], grid[154], grid[155], grid[156], grid[186], grid[188], grid[218], grid[219], grid[220], grid[187]);
evolve8 e188 (grid_evolve[188], grid[155], grid[156], grid[157], grid[187], grid[189], grid[219], grid[220], grid[221], grid[188]);
evolve8 e189 (grid_evolve[189], grid[156], grid[157], grid[158], grid[188], grid[190], grid[220], grid[221], grid[222], grid[189]);
evolve8 e190 (grid_evolve[190], grid[157], grid[158], grid[159], grid[189], grid[191], grid[221], grid[222], grid[223], grid[190]);
evolve5 e191 (grid_evolve[191], grid[158], grid[159], grid[190], grid[222], grid[223], grid[191]);

evolve5 e192 (grid_evolve[192], grid[160], grid[161], grid[193], grid[224], grid[225], grid[192]);
evolve8 e193 (grid_evolve[193], grid[160], grid[161], grid[162], grid[192], grid[194], grid[224], grid[225], grid[226], grid[193]);
evolve8 e194 (grid_evolve[194], grid[161], grid[162], grid[163], grid[193], grid[195], grid[225], grid[226], grid[227], grid[194]);
evolve8 e195 (grid_evolve[195], grid[162], grid[163], grid[164], grid[194], grid[196], grid[226], grid[227], grid[228], grid[195]);
evolve8 e196 (grid_evolve[196], grid[163], grid[164], grid[165], grid[195], grid[197], grid[227], grid[228], grid[229], grid[196]);
evolve8 e197 (grid_evolve[197], grid[164], grid[165], grid[166], grid[196], grid[198], grid[228], grid[229], grid[230], grid[197]);
evolve8 e198 (grid_evolve[198], grid[165], grid[166], grid[167], grid[197], grid[199], grid[229], grid[230], grid[231], grid[198]);
evolve8 e199 (grid_evolve[199], grid[166], grid[167], grid[168], grid[198], grid[200], grid[230], grid[231], grid[232], grid[199]);
evolve8 e200 (grid_evolve[200], grid[167], grid[168], grid[169], grid[199], grid[201], grid[231], grid[232], grid[233], grid[200]);
evolve8 e201 (grid_evolve[201], grid[168], grid[169], grid[170], grid[200], grid[202], grid[232], grid[233], grid[234], grid[201]);
evolve8 e202 (grid_evolve[202], grid[169], grid[170], grid[171], grid[201], grid[203], grid[233], grid[234], grid[235], grid[202]);
evolve8 e203 (grid_evolve[203], grid[170], grid[171], grid[172], grid[202], grid[204], grid[234], grid[235], grid[236], grid[203]);
evolve8 e204 (grid_evolve[204], grid[171], grid[172], grid[173], grid[203], grid[205], grid[235], grid[236], grid[237], grid[204]);
evolve8 e205 (grid_evolve[205], grid[172], grid[173], grid[174], grid[204], grid[206], grid[236], grid[237], grid[238], grid[205]);
evolve8 e206 (grid_evolve[206], grid[173], grid[174], grid[175], grid[205], grid[207], grid[237], grid[238], grid[239], grid[206]);
evolve8 e207 (grid_evolve[207], grid[174], grid[175], grid[176], grid[206], grid[208], grid[238], grid[239], grid[240], grid[207]);
evolve8 e208 (grid_evolve[208], grid[175], grid[176], grid[177], grid[207], grid[209], grid[239], grid[240], grid[241], grid[208]);
evolve8 e209 (grid_evolve[209], grid[176], grid[177], grid[178], grid[208], grid[210], grid[240], grid[241], grid[242], grid[209]);
evolve8 e210 (grid_evolve[210], grid[177], grid[178], grid[179], grid[209], grid[211], grid[241], grid[242], grid[243], grid[210]);
evolve8 e211 (grid_evolve[211], grid[178], grid[179], grid[180], grid[210], grid[212], grid[242], grid[243], grid[244], grid[211]);
evolve8 e212 (grid_evolve[212], grid[179], grid[180], grid[181], grid[211], grid[213], grid[243], grid[244], grid[245], grid[212]);
evolve8 e213 (grid_evolve[213], grid[180], grid[181], grid[182], grid[212], grid[214], grid[244], grid[245], grid[246], grid[213]);
evolve8 e214 (grid_evolve[214], grid[181], grid[182], grid[183], grid[213], grid[215], grid[245], grid[246], grid[247], grid[214]);
evolve8 e215 (grid_evolve[215], grid[182], grid[183], grid[184], grid[214], grid[216], grid[246], grid[247], grid[248], grid[215]);
evolve8 e216 (grid_evolve[216], grid[183], grid[184], grid[185], grid[215], grid[217], grid[247], grid[248], grid[249], grid[216]);
evolve8 e217 (grid_evolve[217], grid[184], grid[185], grid[186], grid[216], grid[218], grid[248], grid[249], grid[250], grid[217]);
evolve8 e218 (grid_evolve[218], grid[185], grid[186], grid[187], grid[217], grid[219], grid[249], grid[250], grid[251], grid[218]);
evolve8 e219 (grid_evolve[219], grid[186], grid[187], grid[188], grid[218], grid[220], grid[250], grid[251], grid[252], grid[219]);
evolve8 e220 (grid_evolve[220], grid[187], grid[188], grid[189], grid[219], grid[221], grid[251], grid[252], grid[253], grid[220]);
evolve8 e221 (grid_evolve[221], grid[188], grid[189], grid[190], grid[220], grid[222], grid[252], grid[253], grid[254], grid[221]);
evolve8 e222 (grid_evolve[222], grid[189], grid[190], grid[191], grid[221], grid[223], grid[253], grid[254], grid[255], grid[222]);
evolve5 e223 (grid_evolve[223], grid[190], grid[191], grid[222], grid[254], grid[255], grid[223]);

evolve5 e224 (grid_evolve[224], grid[192], grid[193], grid[225], grid[256], grid[257], grid[224]);
evolve8 e225 (grid_evolve[225], grid[192], grid[193], grid[194], grid[224], grid[226], grid[256], grid[257], grid[258], grid[225]);
evolve8 e226 (grid_evolve[226], grid[193], grid[194], grid[195], grid[225], grid[227], grid[257], grid[258], grid[259], grid[226]);
evolve8 e227 (grid_evolve[227], grid[194], grid[195], grid[196], grid[226], grid[228], grid[258], grid[259], grid[260], grid[227]);
evolve8 e228 (grid_evolve[228], grid[195], grid[196], grid[197], grid[227], grid[229], grid[259], grid[260], grid[261], grid[228]);
evolve8 e229 (grid_evolve[229], grid[196], grid[197], grid[198], grid[228], grid[230], grid[260], grid[261], grid[262], grid[229]);
evolve8 e230 (grid_evolve[230], grid[197], grid[198], grid[199], grid[229], grid[231], grid[261], grid[262], grid[263], grid[230]);
evolve8 e231 (grid_evolve[231], grid[198], grid[199], grid[200], grid[230], grid[232], grid[262], grid[263], grid[264], grid[231]);
evolve8 e232 (grid_evolve[232], grid[199], grid[200], grid[201], grid[231], grid[233], grid[263], grid[264], grid[265], grid[232]);
evolve8 e233 (grid_evolve[233], grid[200], grid[201], grid[202], grid[232], grid[234], grid[264], grid[265], grid[266], grid[233]);
evolve8 e234 (grid_evolve[234], grid[201], grid[202], grid[203], grid[233], grid[235], grid[265], grid[266], grid[267], grid[234]);
evolve8 e235 (grid_evolve[235], grid[202], grid[203], grid[204], grid[234], grid[236], grid[266], grid[267], grid[268], grid[235]);
evolve8 e236 (grid_evolve[236], grid[203], grid[204], grid[205], grid[235], grid[237], grid[267], grid[268], grid[269], grid[236]);
evolve8 e237 (grid_evolve[237], grid[204], grid[205], grid[206], grid[236], grid[238], grid[268], grid[269], grid[270], grid[237]);
evolve8 e238 (grid_evolve[238], grid[205], grid[206], grid[207], grid[237], grid[239], grid[269], grid[270], grid[271], grid[238]);
evolve8 e239 (grid_evolve[239], grid[206], grid[207], grid[208], grid[238], grid[240], grid[270], grid[271], grid[272], grid[239]);
evolve8 e240 (grid_evolve[240], grid[207], grid[208], grid[209], grid[239], grid[241], grid[271], grid[272], grid[273], grid[240]);
evolve8 e241 (grid_evolve[241], grid[208], grid[209], grid[210], grid[240], grid[242], grid[272], grid[273], grid[274], grid[241]);
evolve8 e242 (grid_evolve[242], grid[209], grid[210], grid[211], grid[241], grid[243], grid[273], grid[274], grid[275], grid[242]);
evolve8 e243 (grid_evolve[243], grid[210], grid[211], grid[212], grid[242], grid[244], grid[274], grid[275], grid[276], grid[243]);
evolve8 e244 (grid_evolve[244], grid[211], grid[212], grid[213], grid[243], grid[245], grid[275], grid[276], grid[277], grid[244]);
evolve8 e245 (grid_evolve[245], grid[212], grid[213], grid[214], grid[244], grid[246], grid[276], grid[277], grid[278], grid[245]);
evolve8 e246 (grid_evolve[246], grid[213], grid[214], grid[215], grid[245], grid[247], grid[277], grid[278], grid[279], grid[246]);
evolve8 e247 (grid_evolve[247], grid[214], grid[215], grid[216], grid[246], grid[248], grid[278], grid[279], grid[280], grid[247]);
evolve8 e248 (grid_evolve[248], grid[215], grid[216], grid[217], grid[247], grid[249], grid[279], grid[280], grid[281], grid[248]);
evolve8 e249 (grid_evolve[249], grid[216], grid[217], grid[218], grid[248], grid[250], grid[280], grid[281], grid[282], grid[249]);
evolve8 e250 (grid_evolve[250], grid[217], grid[218], grid[219], grid[249], grid[251], grid[281], grid[282], grid[283], grid[250]);
evolve8 e251 (grid_evolve[251], grid[218], grid[219], grid[220], grid[250], grid[252], grid[282], grid[283], grid[284], grid[251]);
evolve8 e252 (grid_evolve[252], grid[219], grid[220], grid[221], grid[251], grid[253], grid[283], grid[284], grid[285], grid[252]);
evolve8 e253 (grid_evolve[253], grid[220], grid[221], grid[222], grid[252], grid[254], grid[284], grid[285], grid[286], grid[253]);
evolve8 e254 (grid_evolve[254], grid[221], grid[222], grid[223], grid[253], grid[255], grid[285], grid[286], grid[287], grid[254]);
evolve5 e255 (grid_evolve[255], grid[222], grid[223], grid[254], grid[286], grid[287], grid[255]);

evolve5 e256 (grid_evolve[256], grid[224], grid[225], grid[257], grid[288], grid[289], grid[256]);
evolve8 e257 (grid_evolve[257], grid[224], grid[225], grid[226], grid[256], grid[258], grid[288], grid[289], grid[290], grid[257]);
evolve8 e258 (grid_evolve[258], grid[225], grid[226], grid[227], grid[257], grid[259], grid[289], grid[290], grid[291], grid[258]);
evolve8 e259 (grid_evolve[259], grid[226], grid[227], grid[228], grid[258], grid[260], grid[290], grid[291], grid[292], grid[259]);
evolve8 e260 (grid_evolve[260], grid[227], grid[228], grid[229], grid[259], grid[261], grid[291], grid[292], grid[293], grid[260]);
evolve8 e261 (grid_evolve[261], grid[228], grid[229], grid[230], grid[260], grid[262], grid[292], grid[293], grid[294], grid[261]);
evolve8 e262 (grid_evolve[262], grid[229], grid[230], grid[231], grid[261], grid[263], grid[293], grid[294], grid[295], grid[262]);
evolve8 e263 (grid_evolve[263], grid[230], grid[231], grid[232], grid[262], grid[264], grid[294], grid[295], grid[296], grid[263]);
evolve8 e264 (grid_evolve[264], grid[231], grid[232], grid[233], grid[263], grid[265], grid[295], grid[296], grid[297], grid[264]);
evolve8 e265 (grid_evolve[265], grid[232], grid[233], grid[234], grid[264], grid[266], grid[296], grid[297], grid[298], grid[265]);
evolve8 e266 (grid_evolve[266], grid[233], grid[234], grid[235], grid[265], grid[267], grid[297], grid[298], grid[299], grid[266]);
evolve8 e267 (grid_evolve[267], grid[234], grid[235], grid[236], grid[266], grid[268], grid[298], grid[299], grid[300], grid[267]);
evolve8 e268 (grid_evolve[268], grid[235], grid[236], grid[237], grid[267], grid[269], grid[299], grid[300], grid[301], grid[268]);
evolve8 e269 (grid_evolve[269], grid[236], grid[237], grid[238], grid[268], grid[270], grid[300], grid[301], grid[302], grid[269]);
evolve8 e270 (grid_evolve[270], grid[237], grid[238], grid[239], grid[269], grid[271], grid[301], grid[302], grid[303], grid[270]);
evolve8 e271 (grid_evolve[271], grid[238], grid[239], grid[240], grid[270], grid[272], grid[302], grid[303], grid[304], grid[271]);
evolve8 e272 (grid_evolve[272], grid[239], grid[240], grid[241], grid[271], grid[273], grid[303], grid[304], grid[305], grid[272]);
evolve8 e273 (grid_evolve[273], grid[240], grid[241], grid[242], grid[272], grid[274], grid[304], grid[305], grid[306], grid[273]);
evolve8 e274 (grid_evolve[274], grid[241], grid[242], grid[243], grid[273], grid[275], grid[305], grid[306], grid[307], grid[274]);
evolve8 e275 (grid_evolve[275], grid[242], grid[243], grid[244], grid[274], grid[276], grid[306], grid[307], grid[308], grid[275]);
evolve8 e276 (grid_evolve[276], grid[243], grid[244], grid[245], grid[275], grid[277], grid[307], grid[308], grid[309], grid[276]);
evolve8 e277 (grid_evolve[277], grid[244], grid[245], grid[246], grid[276], grid[278], grid[308], grid[309], grid[310], grid[277]);
evolve8 e278 (grid_evolve[278], grid[245], grid[246], grid[247], grid[277], grid[279], grid[309], grid[310], grid[311], grid[278]);
evolve8 e279 (grid_evolve[279], grid[246], grid[247], grid[248], grid[278], grid[280], grid[310], grid[311], grid[312], grid[279]);
evolve8 e280 (grid_evolve[280], grid[247], grid[248], grid[249], grid[279], grid[281], grid[311], grid[312], grid[313], grid[280]);
evolve8 e281 (grid_evolve[281], grid[248], grid[249], grid[250], grid[280], grid[282], grid[312], grid[313], grid[314], grid[281]);
evolve8 e282 (grid_evolve[282], grid[249], grid[250], grid[251], grid[281], grid[283], grid[313], grid[314], grid[315], grid[282]);
evolve8 e283 (grid_evolve[283], grid[250], grid[251], grid[252], grid[282], grid[284], grid[314], grid[315], grid[316], grid[283]);
evolve8 e284 (grid_evolve[284], grid[251], grid[252], grid[253], grid[283], grid[285], grid[315], grid[316], grid[317], grid[284]);
evolve8 e285 (grid_evolve[285], grid[252], grid[253], grid[254], grid[284], grid[286], grid[316], grid[317], grid[318], grid[285]);
evolve8 e286 (grid_evolve[286], grid[253], grid[254], grid[255], grid[285], grid[287], grid[317], grid[318], grid[319], grid[286]);
evolve5 e287 (grid_evolve[287], grid[254], grid[255], grid[286], grid[318], grid[319], grid[287]);

evolve5 e288 (grid_evolve[288], grid[256], grid[257], grid[289], grid[320], grid[321], grid[288]);
evolve8 e289 (grid_evolve[289], grid[256], grid[257], grid[258], grid[288], grid[290], grid[320], grid[321], grid[322], grid[289]);
evolve8 e290 (grid_evolve[290], grid[257], grid[258], grid[259], grid[289], grid[291], grid[321], grid[322], grid[323], grid[290]);
evolve8 e291 (grid_evolve[291], grid[258], grid[259], grid[260], grid[290], grid[292], grid[322], grid[323], grid[324], grid[291]);
evolve8 e292 (grid_evolve[292], grid[259], grid[260], grid[261], grid[291], grid[293], grid[323], grid[324], grid[325], grid[292]);
evolve8 e293 (grid_evolve[293], grid[260], grid[261], grid[262], grid[292], grid[294], grid[324], grid[325], grid[326], grid[293]);
evolve8 e294 (grid_evolve[294], grid[261], grid[262], grid[263], grid[293], grid[295], grid[325], grid[326], grid[327], grid[294]);
evolve8 e295 (grid_evolve[295], grid[262], grid[263], grid[264], grid[294], grid[296], grid[326], grid[327], grid[328], grid[295]);
evolve8 e296 (grid_evolve[296], grid[263], grid[264], grid[265], grid[295], grid[297], grid[327], grid[328], grid[329], grid[296]);
evolve8 e297 (grid_evolve[297], grid[264], grid[265], grid[266], grid[296], grid[298], grid[328], grid[329], grid[330], grid[297]);
evolve8 e298 (grid_evolve[298], grid[265], grid[266], grid[267], grid[297], grid[299], grid[329], grid[330], grid[331], grid[298]);
evolve8 e299 (grid_evolve[299], grid[266], grid[267], grid[268], grid[298], grid[300], grid[330], grid[331], grid[332], grid[299]);
evolve8 e300 (grid_evolve[300], grid[267], grid[268], grid[269], grid[299], grid[301], grid[331], grid[332], grid[333], grid[300]);
evolve8 e301 (grid_evolve[301], grid[268], grid[269], grid[270], grid[300], grid[302], grid[332], grid[333], grid[334], grid[301]);
evolve8 e302 (grid_evolve[302], grid[269], grid[270], grid[271], grid[301], grid[303], grid[333], grid[334], grid[335], grid[302]);
evolve8 e303 (grid_evolve[303], grid[270], grid[271], grid[272], grid[302], grid[304], grid[334], grid[335], grid[336], grid[303]);
evolve8 e304 (grid_evolve[304], grid[271], grid[272], grid[273], grid[303], grid[305], grid[335], grid[336], grid[337], grid[304]);
evolve8 e305 (grid_evolve[305], grid[272], grid[273], grid[274], grid[304], grid[306], grid[336], grid[337], grid[338], grid[305]);
evolve8 e306 (grid_evolve[306], grid[273], grid[274], grid[275], grid[305], grid[307], grid[337], grid[338], grid[339], grid[306]);
evolve8 e307 (grid_evolve[307], grid[274], grid[275], grid[276], grid[306], grid[308], grid[338], grid[339], grid[340], grid[307]);
evolve8 e308 (grid_evolve[308], grid[275], grid[276], grid[277], grid[307], grid[309], grid[339], grid[340], grid[341], grid[308]);
evolve8 e309 (grid_evolve[309], grid[276], grid[277], grid[278], grid[308], grid[310], grid[340], grid[341], grid[342], grid[309]);
evolve8 e310 (grid_evolve[310], grid[277], grid[278], grid[279], grid[309], grid[311], grid[341], grid[342], grid[343], grid[310]);
evolve8 e311 (grid_evolve[311], grid[278], grid[279], grid[280], grid[310], grid[312], grid[342], grid[343], grid[344], grid[311]);
evolve8 e312 (grid_evolve[312], grid[279], grid[280], grid[281], grid[311], grid[313], grid[343], grid[344], grid[345], grid[312]);
evolve8 e313 (grid_evolve[313], grid[280], grid[281], grid[282], grid[312], grid[314], grid[344], grid[345], grid[346], grid[313]);
evolve8 e314 (grid_evolve[314], grid[281], grid[282], grid[283], grid[313], grid[315], grid[345], grid[346], grid[347], grid[314]);
evolve8 e315 (grid_evolve[315], grid[282], grid[283], grid[284], grid[314], grid[316], grid[346], grid[347], grid[348], grid[315]);
evolve8 e316 (grid_evolve[316], grid[283], grid[284], grid[285], grid[315], grid[317], grid[347], grid[348], grid[349], grid[316]);
evolve8 e317 (grid_evolve[317], grid[284], grid[285], grid[286], grid[316], grid[318], grid[348], grid[349], grid[350], grid[317]);
evolve8 e318 (grid_evolve[318], grid[285], grid[286], grid[287], grid[317], grid[319], grid[349], grid[350], grid[351], grid[318]);
evolve5 e319 (grid_evolve[319], grid[286], grid[287], grid[318], grid[350], grid[351], grid[319]);

evolve5 e320 (grid_evolve[320], grid[288], grid[289], grid[321], grid[352], grid[353], grid[320]);
evolve8 e321 (grid_evolve[321], grid[288], grid[289], grid[290], grid[320], grid[322], grid[352], grid[353], grid[354], grid[321]);
evolve8 e322 (grid_evolve[322], grid[289], grid[290], grid[291], grid[321], grid[323], grid[353], grid[354], grid[355], grid[322]);
evolve8 e323 (grid_evolve[323], grid[290], grid[291], grid[292], grid[322], grid[324], grid[354], grid[355], grid[356], grid[323]);
evolve8 e324 (grid_evolve[324], grid[291], grid[292], grid[293], grid[323], grid[325], grid[355], grid[356], grid[357], grid[324]);
evolve8 e325 (grid_evolve[325], grid[292], grid[293], grid[294], grid[324], grid[326], grid[356], grid[357], grid[358], grid[325]);
evolve8 e326 (grid_evolve[326], grid[293], grid[294], grid[295], grid[325], grid[327], grid[357], grid[358], grid[359], grid[326]);
evolve8 e327 (grid_evolve[327], grid[294], grid[295], grid[296], grid[326], grid[328], grid[358], grid[359], grid[360], grid[327]);
evolve8 e328 (grid_evolve[328], grid[295], grid[296], grid[297], grid[327], grid[329], grid[359], grid[360], grid[361], grid[328]);
evolve8 e329 (grid_evolve[329], grid[296], grid[297], grid[298], grid[328], grid[330], grid[360], grid[361], grid[362], grid[329]);
evolve8 e330 (grid_evolve[330], grid[297], grid[298], grid[299], grid[329], grid[331], grid[361], grid[362], grid[363], grid[330]);
evolve8 e331 (grid_evolve[331], grid[298], grid[299], grid[300], grid[330], grid[332], grid[362], grid[363], grid[364], grid[331]);
evolve8 e332 (grid_evolve[332], grid[299], grid[300], grid[301], grid[331], grid[333], grid[363], grid[364], grid[365], grid[332]);
evolve8 e333 (grid_evolve[333], grid[300], grid[301], grid[302], grid[332], grid[334], grid[364], grid[365], grid[366], grid[333]);
evolve8 e334 (grid_evolve[334], grid[301], grid[302], grid[303], grid[333], grid[335], grid[365], grid[366], grid[367], grid[334]);
evolve8 e335 (grid_evolve[335], grid[302], grid[303], grid[304], grid[334], grid[336], grid[366], grid[367], grid[368], grid[335]);
evolve8 e336 (grid_evolve[336], grid[303], grid[304], grid[305], grid[335], grid[337], grid[367], grid[368], grid[369], grid[336]);
evolve8 e337 (grid_evolve[337], grid[304], grid[305], grid[306], grid[336], grid[338], grid[368], grid[369], grid[370], grid[337]);
evolve8 e338 (grid_evolve[338], grid[305], grid[306], grid[307], grid[337], grid[339], grid[369], grid[370], grid[371], grid[338]);
evolve8 e339 (grid_evolve[339], grid[306], grid[307], grid[308], grid[338], grid[340], grid[370], grid[371], grid[372], grid[339]);
evolve8 e340 (grid_evolve[340], grid[307], grid[308], grid[309], grid[339], grid[341], grid[371], grid[372], grid[373], grid[340]);
evolve8 e341 (grid_evolve[341], grid[308], grid[309], grid[310], grid[340], grid[342], grid[372], grid[373], grid[374], grid[341]);
evolve8 e342 (grid_evolve[342], grid[309], grid[310], grid[311], grid[341], grid[343], grid[373], grid[374], grid[375], grid[342]);
evolve8 e343 (grid_evolve[343], grid[310], grid[311], grid[312], grid[342], grid[344], grid[374], grid[375], grid[376], grid[343]);
evolve8 e344 (grid_evolve[344], grid[311], grid[312], grid[313], grid[343], grid[345], grid[375], grid[376], grid[377], grid[344]);
evolve8 e345 (grid_evolve[345], grid[312], grid[313], grid[314], grid[344], grid[346], grid[376], grid[377], grid[378], grid[345]);
evolve8 e346 (grid_evolve[346], grid[313], grid[314], grid[315], grid[345], grid[347], grid[377], grid[378], grid[379], grid[346]);
evolve8 e347 (grid_evolve[347], grid[314], grid[315], grid[316], grid[346], grid[348], grid[378], grid[379], grid[380], grid[347]);
evolve8 e348 (grid_evolve[348], grid[315], grid[316], grid[317], grid[347], grid[349], grid[379], grid[380], grid[381], grid[348]);
evolve8 e349 (grid_evolve[349], grid[316], grid[317], grid[318], grid[348], grid[350], grid[380], grid[381], grid[382], grid[349]);
evolve8 e350 (grid_evolve[350], grid[317], grid[318], grid[319], grid[349], grid[351], grid[381], grid[382], grid[383], grid[350]);
evolve5 e351 (grid_evolve[351], grid[318], grid[319], grid[350], grid[382], grid[383], grid[351]);

evolve5 e352 (grid_evolve[352], grid[320], grid[321], grid[353], grid[384], grid[385], grid[352]);
evolve8 e353 (grid_evolve[353], grid[320], grid[321], grid[322], grid[352], grid[354], grid[384], grid[385], grid[386], grid[353]);
evolve8 e354 (grid_evolve[354], grid[321], grid[322], grid[323], grid[353], grid[355], grid[385], grid[386], grid[387], grid[354]);
evolve8 e355 (grid_evolve[355], grid[322], grid[323], grid[324], grid[354], grid[356], grid[386], grid[387], grid[388], grid[355]);
evolve8 e356 (grid_evolve[356], grid[323], grid[324], grid[325], grid[355], grid[357], grid[387], grid[388], grid[389], grid[356]);
evolve8 e357 (grid_evolve[357], grid[324], grid[325], grid[326], grid[356], grid[358], grid[388], grid[389], grid[390], grid[357]);
evolve8 e358 (grid_evolve[358], grid[325], grid[326], grid[327], grid[357], grid[359], grid[389], grid[390], grid[391], grid[358]);
evolve8 e359 (grid_evolve[359], grid[326], grid[327], grid[328], grid[358], grid[360], grid[390], grid[391], grid[392], grid[359]);
evolve8 e360 (grid_evolve[360], grid[327], grid[328], grid[329], grid[359], grid[361], grid[391], grid[392], grid[393], grid[360]);
evolve8 e361 (grid_evolve[361], grid[328], grid[329], grid[330], grid[360], grid[362], grid[392], grid[393], grid[394], grid[361]);
evolve8 e362 (grid_evolve[362], grid[329], grid[330], grid[331], grid[361], grid[363], grid[393], grid[394], grid[395], grid[362]);
evolve8 e363 (grid_evolve[363], grid[330], grid[331], grid[332], grid[362], grid[364], grid[394], grid[395], grid[396], grid[363]);
evolve8 e364 (grid_evolve[364], grid[331], grid[332], grid[333], grid[363], grid[365], grid[395], grid[396], grid[397], grid[364]);
evolve8 e365 (grid_evolve[365], grid[332], grid[333], grid[334], grid[364], grid[366], grid[396], grid[397], grid[398], grid[365]);
evolve8 e366 (grid_evolve[366], grid[333], grid[334], grid[335], grid[365], grid[367], grid[397], grid[398], grid[399], grid[366]);
evolve8 e367 (grid_evolve[367], grid[334], grid[335], grid[336], grid[366], grid[368], grid[398], grid[399], grid[400], grid[367]);
evolve8 e368 (grid_evolve[368], grid[335], grid[336], grid[337], grid[367], grid[369], grid[399], grid[400], grid[401], grid[368]);
evolve8 e369 (grid_evolve[369], grid[336], grid[337], grid[338], grid[368], grid[370], grid[400], grid[401], grid[402], grid[369]);
evolve8 e370 (grid_evolve[370], grid[337], grid[338], grid[339], grid[369], grid[371], grid[401], grid[402], grid[403], grid[370]);
evolve8 e371 (grid_evolve[371], grid[338], grid[339], grid[340], grid[370], grid[372], grid[402], grid[403], grid[404], grid[371]);
evolve8 e372 (grid_evolve[372], grid[339], grid[340], grid[341], grid[371], grid[373], grid[403], grid[404], grid[405], grid[372]);
evolve8 e373 (grid_evolve[373], grid[340], grid[341], grid[342], grid[372], grid[374], grid[404], grid[405], grid[406], grid[373]);
evolve8 e374 (grid_evolve[374], grid[341], grid[342], grid[343], grid[373], grid[375], grid[405], grid[406], grid[407], grid[374]);
evolve8 e375 (grid_evolve[375], grid[342], grid[343], grid[344], grid[374], grid[376], grid[406], grid[407], grid[408], grid[375]);
evolve8 e376 (grid_evolve[376], grid[343], grid[344], grid[345], grid[375], grid[377], grid[407], grid[408], grid[409], grid[376]);
evolve8 e377 (grid_evolve[377], grid[344], grid[345], grid[346], grid[376], grid[378], grid[408], grid[409], grid[410], grid[377]);
evolve8 e378 (grid_evolve[378], grid[345], grid[346], grid[347], grid[377], grid[379], grid[409], grid[410], grid[411], grid[378]);
evolve8 e379 (grid_evolve[379], grid[346], grid[347], grid[348], grid[378], grid[380], grid[410], grid[411], grid[412], grid[379]);
evolve8 e380 (grid_evolve[380], grid[347], grid[348], grid[349], grid[379], grid[381], grid[411], grid[412], grid[413], grid[380]);
evolve8 e381 (grid_evolve[381], grid[348], grid[349], grid[350], grid[380], grid[382], grid[412], grid[413], grid[414], grid[381]);
evolve8 e382 (grid_evolve[382], grid[349], grid[350], grid[351], grid[381], grid[383], grid[413], grid[414], grid[415], grid[382]);
evolve5 e383 (grid_evolve[383], grid[350], grid[351], grid[382], grid[414], grid[415], grid[383]);

evolve5 e384 (grid_evolve[384], grid[352], grid[353], grid[385], grid[416], grid[417], grid[384]);
evolve8 e385 (grid_evolve[385], grid[352], grid[353], grid[354], grid[384], grid[386], grid[416], grid[417], grid[418], grid[385]);
evolve8 e386 (grid_evolve[386], grid[353], grid[354], grid[355], grid[385], grid[387], grid[417], grid[418], grid[419], grid[386]);
evolve8 e387 (grid_evolve[387], grid[354], grid[355], grid[356], grid[386], grid[388], grid[418], grid[419], grid[420], grid[387]);
evolve8 e388 (grid_evolve[388], grid[355], grid[356], grid[357], grid[387], grid[389], grid[419], grid[420], grid[421], grid[388]);
evolve8 e389 (grid_evolve[389], grid[356], grid[357], grid[358], grid[388], grid[390], grid[420], grid[421], grid[422], grid[389]);
evolve8 e390 (grid_evolve[390], grid[357], grid[358], grid[359], grid[389], grid[391], grid[421], grid[422], grid[423], grid[390]);
evolve8 e391 (grid_evolve[391], grid[358], grid[359], grid[360], grid[390], grid[392], grid[422], grid[423], grid[424], grid[391]);
evolve8 e392 (grid_evolve[392], grid[359], grid[360], grid[361], grid[391], grid[393], grid[423], grid[424], grid[425], grid[392]);
evolve8 e393 (grid_evolve[393], grid[360], grid[361], grid[362], grid[392], grid[394], grid[424], grid[425], grid[426], grid[393]);
evolve8 e394 (grid_evolve[394], grid[361], grid[362], grid[363], grid[393], grid[395], grid[425], grid[426], grid[427], grid[394]);
evolve8 e395 (grid_evolve[395], grid[362], grid[363], grid[364], grid[394], grid[396], grid[426], grid[427], grid[428], grid[395]);
evolve8 e396 (grid_evolve[396], grid[363], grid[364], grid[365], grid[395], grid[397], grid[427], grid[428], grid[429], grid[396]);
evolve8 e397 (grid_evolve[397], grid[364], grid[365], grid[366], grid[396], grid[398], grid[428], grid[429], grid[430], grid[397]);
evolve8 e398 (grid_evolve[398], grid[365], grid[366], grid[367], grid[397], grid[399], grid[429], grid[430], grid[431], grid[398]);
evolve8 e399 (grid_evolve[399], grid[366], grid[367], grid[368], grid[398], grid[400], grid[430], grid[431], grid[432], grid[399]);
evolve8 e400 (grid_evolve[400], grid[367], grid[368], grid[369], grid[399], grid[401], grid[431], grid[432], grid[433], grid[400]);
evolve8 e401 (grid_evolve[401], grid[368], grid[369], grid[370], grid[400], grid[402], grid[432], grid[433], grid[434], grid[401]);
evolve8 e402 (grid_evolve[402], grid[369], grid[370], grid[371], grid[401], grid[403], grid[433], grid[434], grid[435], grid[402]);
evolve8 e403 (grid_evolve[403], grid[370], grid[371], grid[372], grid[402], grid[404], grid[434], grid[435], grid[436], grid[403]);
evolve8 e404 (grid_evolve[404], grid[371], grid[372], grid[373], grid[403], grid[405], grid[435], grid[436], grid[437], grid[404]);
evolve8 e405 (grid_evolve[405], grid[372], grid[373], grid[374], grid[404], grid[406], grid[436], grid[437], grid[438], grid[405]);
evolve8 e406 (grid_evolve[406], grid[373], grid[374], grid[375], grid[405], grid[407], grid[437], grid[438], grid[439], grid[406]);
evolve8 e407 (grid_evolve[407], grid[374], grid[375], grid[376], grid[406], grid[408], grid[438], grid[439], grid[440], grid[407]);
evolve8 e408 (grid_evolve[408], grid[375], grid[376], grid[377], grid[407], grid[409], grid[439], grid[440], grid[441], grid[408]);
evolve8 e409 (grid_evolve[409], grid[376], grid[377], grid[378], grid[408], grid[410], grid[440], grid[441], grid[442], grid[409]);
evolve8 e410 (grid_evolve[410], grid[377], grid[378], grid[379], grid[409], grid[411], grid[441], grid[442], grid[443], grid[410]);
evolve8 e411 (grid_evolve[411], grid[378], grid[379], grid[380], grid[410], grid[412], grid[442], grid[443], grid[444], grid[411]);
evolve8 e412 (grid_evolve[412], grid[379], grid[380], grid[381], grid[411], grid[413], grid[443], grid[444], grid[445], grid[412]);
evolve8 e413 (grid_evolve[413], grid[380], grid[381], grid[382], grid[412], grid[414], grid[444], grid[445], grid[446], grid[413]);
evolve8 e414 (grid_evolve[414], grid[381], grid[382], grid[383], grid[413], grid[415], grid[445], grid[446], grid[447], grid[414]);
evolve5 e415 (grid_evolve[415], grid[382], grid[383], grid[414], grid[446], grid[447], grid[415]);

evolve5 e416 (grid_evolve[416], grid[384], grid[385], grid[417], grid[448], grid[449], grid[416]);
evolve8 e417 (grid_evolve[417], grid[384], grid[385], grid[386], grid[416], grid[418], grid[448], grid[449], grid[450], grid[417]);
evolve8 e418 (grid_evolve[418], grid[385], grid[386], grid[387], grid[417], grid[419], grid[449], grid[450], grid[451], grid[418]);
evolve8 e419 (grid_evolve[419], grid[386], grid[387], grid[388], grid[418], grid[420], grid[450], grid[451], grid[452], grid[419]);
evolve8 e420 (grid_evolve[420], grid[387], grid[388], grid[389], grid[419], grid[421], grid[451], grid[452], grid[453], grid[420]);
evolve8 e421 (grid_evolve[421], grid[388], grid[389], grid[390], grid[420], grid[422], grid[452], grid[453], grid[454], grid[421]);
evolve8 e422 (grid_evolve[422], grid[389], grid[390], grid[391], grid[421], grid[423], grid[453], grid[454], grid[455], grid[422]);
evolve8 e423 (grid_evolve[423], grid[390], grid[391], grid[392], grid[422], grid[424], grid[454], grid[455], grid[456], grid[423]);
evolve8 e424 (grid_evolve[424], grid[391], grid[392], grid[393], grid[423], grid[425], grid[455], grid[456], grid[457], grid[424]);
evolve8 e425 (grid_evolve[425], grid[392], grid[393], grid[394], grid[424], grid[426], grid[456], grid[457], grid[458], grid[425]);
evolve8 e426 (grid_evolve[426], grid[393], grid[394], grid[395], grid[425], grid[427], grid[457], grid[458], grid[459], grid[426]);
evolve8 e427 (grid_evolve[427], grid[394], grid[395], grid[396], grid[426], grid[428], grid[458], grid[459], grid[460], grid[427]);
evolve8 e428 (grid_evolve[428], grid[395], grid[396], grid[397], grid[427], grid[429], grid[459], grid[460], grid[461], grid[428]);
evolve8 e429 (grid_evolve[429], grid[396], grid[397], grid[398], grid[428], grid[430], grid[460], grid[461], grid[462], grid[429]);
evolve8 e430 (grid_evolve[430], grid[397], grid[398], grid[399], grid[429], grid[431], grid[461], grid[462], grid[463], grid[430]);
evolve8 e431 (grid_evolve[431], grid[398], grid[399], grid[400], grid[430], grid[432], grid[462], grid[463], grid[464], grid[431]);
evolve8 e432 (grid_evolve[432], grid[399], grid[400], grid[401], grid[431], grid[433], grid[463], grid[464], grid[465], grid[432]);
evolve8 e433 (grid_evolve[433], grid[400], grid[401], grid[402], grid[432], grid[434], grid[464], grid[465], grid[466], grid[433]);
evolve8 e434 (grid_evolve[434], grid[401], grid[402], grid[403], grid[433], grid[435], grid[465], grid[466], grid[467], grid[434]);
evolve8 e435 (grid_evolve[435], grid[402], grid[403], grid[404], grid[434], grid[436], grid[466], grid[467], grid[468], grid[435]);
evolve8 e436 (grid_evolve[436], grid[403], grid[404], grid[405], grid[435], grid[437], grid[467], grid[468], grid[469], grid[436]);
evolve8 e437 (grid_evolve[437], grid[404], grid[405], grid[406], grid[436], grid[438], grid[468], grid[469], grid[470], grid[437]);
evolve8 e438 (grid_evolve[438], grid[405], grid[406], grid[407], grid[437], grid[439], grid[469], grid[470], grid[471], grid[438]);
evolve8 e439 (grid_evolve[439], grid[406], grid[407], grid[408], grid[438], grid[440], grid[470], grid[471], grid[472], grid[439]);
evolve8 e440 (grid_evolve[440], grid[407], grid[408], grid[409], grid[439], grid[441], grid[471], grid[472], grid[473], grid[440]);
evolve8 e441 (grid_evolve[441], grid[408], grid[409], grid[410], grid[440], grid[442], grid[472], grid[473], grid[474], grid[441]);
evolve8 e442 (grid_evolve[442], grid[409], grid[410], grid[411], grid[441], grid[443], grid[473], grid[474], grid[475], grid[442]);
evolve8 e443 (grid_evolve[443], grid[410], grid[411], grid[412], grid[442], grid[444], grid[474], grid[475], grid[476], grid[443]);
evolve8 e444 (grid_evolve[444], grid[411], grid[412], grid[413], grid[443], grid[445], grid[475], grid[476], grid[477], grid[444]);
evolve8 e445 (grid_evolve[445], grid[412], grid[413], grid[414], grid[444], grid[446], grid[476], grid[477], grid[478], grid[445]);
evolve8 e446 (grid_evolve[446], grid[413], grid[414], grid[415], grid[445], grid[447], grid[477], grid[478], grid[479], grid[446]);
evolve5 e447 (grid_evolve[447], grid[414], grid[415], grid[446], grid[478], grid[479], grid[447]);

evolve5 e448 (grid_evolve[448], grid[416], grid[417], grid[449], grid[480], grid[481], grid[448]);
evolve8 e449 (grid_evolve[449], grid[416], grid[417], grid[418], grid[448], grid[450], grid[480], grid[481], grid[482], grid[449]);
evolve8 e450 (grid_evolve[450], grid[417], grid[418], grid[419], grid[449], grid[451], grid[481], grid[482], grid[483], grid[450]);
evolve8 e451 (grid_evolve[451], grid[418], grid[419], grid[420], grid[450], grid[452], grid[482], grid[483], grid[484], grid[451]);
evolve8 e452 (grid_evolve[452], grid[419], grid[420], grid[421], grid[451], grid[453], grid[483], grid[484], grid[485], grid[452]);
evolve8 e453 (grid_evolve[453], grid[420], grid[421], grid[422], grid[452], grid[454], grid[484], grid[485], grid[486], grid[453]);
evolve8 e454 (grid_evolve[454], grid[421], grid[422], grid[423], grid[453], grid[455], grid[485], grid[486], grid[487], grid[454]);
evolve8 e455 (grid_evolve[455], grid[422], grid[423], grid[424], grid[454], grid[456], grid[486], grid[487], grid[488], grid[455]);
evolve8 e456 (grid_evolve[456], grid[423], grid[424], grid[425], grid[455], grid[457], grid[487], grid[488], grid[489], grid[456]);
evolve8 e457 (grid_evolve[457], grid[424], grid[425], grid[426], grid[456], grid[458], grid[488], grid[489], grid[490], grid[457]);
evolve8 e458 (grid_evolve[458], grid[425], grid[426], grid[427], grid[457], grid[459], grid[489], grid[490], grid[491], grid[458]);
evolve8 e459 (grid_evolve[459], grid[426], grid[427], grid[428], grid[458], grid[460], grid[490], grid[491], grid[492], grid[459]);
evolve8 e460 (grid_evolve[460], grid[427], grid[428], grid[429], grid[459], grid[461], grid[491], grid[492], grid[493], grid[460]);
evolve8 e461 (grid_evolve[461], grid[428], grid[429], grid[430], grid[460], grid[462], grid[492], grid[493], grid[494], grid[461]);
evolve8 e462 (grid_evolve[462], grid[429], grid[430], grid[431], grid[461], grid[463], grid[493], grid[494], grid[495], grid[462]);
evolve8 e463 (grid_evolve[463], grid[430], grid[431], grid[432], grid[462], grid[464], grid[494], grid[495], grid[496], grid[463]);
evolve8 e464 (grid_evolve[464], grid[431], grid[432], grid[433], grid[463], grid[465], grid[495], grid[496], grid[497], grid[464]);
evolve8 e465 (grid_evolve[465], grid[432], grid[433], grid[434], grid[464], grid[466], grid[496], grid[497], grid[498], grid[465]);
evolve8 e466 (grid_evolve[466], grid[433], grid[434], grid[435], grid[465], grid[467], grid[497], grid[498], grid[499], grid[466]);
evolve8 e467 (grid_evolve[467], grid[434], grid[435], grid[436], grid[466], grid[468], grid[498], grid[499], grid[500], grid[467]);
evolve8 e468 (grid_evolve[468], grid[435], grid[436], grid[437], grid[467], grid[469], grid[499], grid[500], grid[501], grid[468]);
evolve8 e469 (grid_evolve[469], grid[436], grid[437], grid[438], grid[468], grid[470], grid[500], grid[501], grid[502], grid[469]);
evolve8 e470 (grid_evolve[470], grid[437], grid[438], grid[439], grid[469], grid[471], grid[501], grid[502], grid[503], grid[470]);
evolve8 e471 (grid_evolve[471], grid[438], grid[439], grid[440], grid[470], grid[472], grid[502], grid[503], grid[504], grid[471]);
evolve8 e472 (grid_evolve[472], grid[439], grid[440], grid[441], grid[471], grid[473], grid[503], grid[504], grid[505], grid[472]);
evolve8 e473 (grid_evolve[473], grid[440], grid[441], grid[442], grid[472], grid[474], grid[504], grid[505], grid[506], grid[473]);
evolve8 e474 (grid_evolve[474], grid[441], grid[442], grid[443], grid[473], grid[475], grid[505], grid[506], grid[507], grid[474]);
evolve8 e475 (grid_evolve[475], grid[442], grid[443], grid[444], grid[474], grid[476], grid[506], grid[507], grid[508], grid[475]);
evolve8 e476 (grid_evolve[476], grid[443], grid[444], grid[445], grid[475], grid[477], grid[507], grid[508], grid[509], grid[476]);
evolve8 e477 (grid_evolve[477], grid[444], grid[445], grid[446], grid[476], grid[478], grid[508], grid[509], grid[510], grid[477]);
evolve8 e478 (grid_evolve[478], grid[445], grid[446], grid[447], grid[477], grid[479], grid[509], grid[510], grid[511], grid[478]);
evolve5 e479 (grid_evolve[479], grid[446], grid[447], grid[478], grid[510], grid[511], grid[479]);

evolve5 e480 (grid_evolve[480], grid[448], grid[449], grid[481], grid[512], grid[513], grid[480]);
evolve8 e481 (grid_evolve[481], grid[448], grid[449], grid[450], grid[480], grid[482], grid[512], grid[513], grid[514], grid[481]);
evolve8 e482 (grid_evolve[482], grid[449], grid[450], grid[451], grid[481], grid[483], grid[513], grid[514], grid[515], grid[482]);
evolve8 e483 (grid_evolve[483], grid[450], grid[451], grid[452], grid[482], grid[484], grid[514], grid[515], grid[516], grid[483]);
evolve8 e484 (grid_evolve[484], grid[451], grid[452], grid[453], grid[483], grid[485], grid[515], grid[516], grid[517], grid[484]);
evolve8 e485 (grid_evolve[485], grid[452], grid[453], grid[454], grid[484], grid[486], grid[516], grid[517], grid[518], grid[485]);
evolve8 e486 (grid_evolve[486], grid[453], grid[454], grid[455], grid[485], grid[487], grid[517], grid[518], grid[519], grid[486]);
evolve8 e487 (grid_evolve[487], grid[454], grid[455], grid[456], grid[486], grid[488], grid[518], grid[519], grid[520], grid[487]);
evolve8 e488 (grid_evolve[488], grid[455], grid[456], grid[457], grid[487], grid[489], grid[519], grid[520], grid[521], grid[488]);
evolve8 e489 (grid_evolve[489], grid[456], grid[457], grid[458], grid[488], grid[490], grid[520], grid[521], grid[522], grid[489]);
evolve8 e490 (grid_evolve[490], grid[457], grid[458], grid[459], grid[489], grid[491], grid[521], grid[522], grid[523], grid[490]);
evolve8 e491 (grid_evolve[491], grid[458], grid[459], grid[460], grid[490], grid[492], grid[522], grid[523], grid[524], grid[491]);
evolve8 e492 (grid_evolve[492], grid[459], grid[460], grid[461], grid[491], grid[493], grid[523], grid[524], grid[525], grid[492]);
evolve8 e493 (grid_evolve[493], grid[460], grid[461], grid[462], grid[492], grid[494], grid[524], grid[525], grid[526], grid[493]);
evolve8 e494 (grid_evolve[494], grid[461], grid[462], grid[463], grid[493], grid[495], grid[525], grid[526], grid[527], grid[494]);
evolve8 e495 (grid_evolve[495], grid[462], grid[463], grid[464], grid[494], grid[496], grid[526], grid[527], grid[528], grid[495]);
evolve8 e496 (grid_evolve[496], grid[463], grid[464], grid[465], grid[495], grid[497], grid[527], grid[528], grid[529], grid[496]);
evolve8 e497 (grid_evolve[497], grid[464], grid[465], grid[466], grid[496], grid[498], grid[528], grid[529], grid[530], grid[497]);
evolve8 e498 (grid_evolve[498], grid[465], grid[466], grid[467], grid[497], grid[499], grid[529], grid[530], grid[531], grid[498]);
evolve8 e499 (grid_evolve[499], grid[466], grid[467], grid[468], grid[498], grid[500], grid[530], grid[531], grid[532], grid[499]);
evolve8 e500 (grid_evolve[500], grid[467], grid[468], grid[469], grid[499], grid[501], grid[531], grid[532], grid[533], grid[500]);
evolve8 e501 (grid_evolve[501], grid[468], grid[469], grid[470], grid[500], grid[502], grid[532], grid[533], grid[534], grid[501]);
evolve8 e502 (grid_evolve[502], grid[469], grid[470], grid[471], grid[501], grid[503], grid[533], grid[534], grid[535], grid[502]);
evolve8 e503 (grid_evolve[503], grid[470], grid[471], grid[472], grid[502], grid[504], grid[534], grid[535], grid[536], grid[503]);
evolve8 e504 (grid_evolve[504], grid[471], grid[472], grid[473], grid[503], grid[505], grid[535], grid[536], grid[537], grid[504]);
evolve8 e505 (grid_evolve[505], grid[472], grid[473], grid[474], grid[504], grid[506], grid[536], grid[537], grid[538], grid[505]);
evolve8 e506 (grid_evolve[506], grid[473], grid[474], grid[475], grid[505], grid[507], grid[537], grid[538], grid[539], grid[506]);
evolve8 e507 (grid_evolve[507], grid[474], grid[475], grid[476], grid[506], grid[508], grid[538], grid[539], grid[540], grid[507]);
evolve8 e508 (grid_evolve[508], grid[475], grid[476], grid[477], grid[507], grid[509], grid[539], grid[540], grid[541], grid[508]);
evolve8 e509 (grid_evolve[509], grid[476], grid[477], grid[478], grid[508], grid[510], grid[540], grid[541], grid[542], grid[509]);
evolve8 e510 (grid_evolve[510], grid[477], grid[478], grid[479], grid[509], grid[511], grid[541], grid[542], grid[543], grid[510]);
evolve5 e511 (grid_evolve[511], grid[478], grid[479], grid[510], grid[542], grid[543], grid[511]);

evolve5 e512 (grid_evolve[512], grid[480], grid[481], grid[513], grid[544], grid[545], grid[512]);
evolve8 e513 (grid_evolve[513], grid[480], grid[481], grid[482], grid[512], grid[514], grid[544], grid[545], grid[546], grid[513]);
evolve8 e514 (grid_evolve[514], grid[481], grid[482], grid[483], grid[513], grid[515], grid[545], grid[546], grid[547], grid[514]);
evolve8 e515 (grid_evolve[515], grid[482], grid[483], grid[484], grid[514], grid[516], grid[546], grid[547], grid[548], grid[515]);
evolve8 e516 (grid_evolve[516], grid[483], grid[484], grid[485], grid[515], grid[517], grid[547], grid[548], grid[549], grid[516]);
evolve8 e517 (grid_evolve[517], grid[484], grid[485], grid[486], grid[516], grid[518], grid[548], grid[549], grid[550], grid[517]);
evolve8 e518 (grid_evolve[518], grid[485], grid[486], grid[487], grid[517], grid[519], grid[549], grid[550], grid[551], grid[518]);
evolve8 e519 (grid_evolve[519], grid[486], grid[487], grid[488], grid[518], grid[520], grid[550], grid[551], grid[552], grid[519]);
evolve8 e520 (grid_evolve[520], grid[487], grid[488], grid[489], grid[519], grid[521], grid[551], grid[552], grid[553], grid[520]);
evolve8 e521 (grid_evolve[521], grid[488], grid[489], grid[490], grid[520], grid[522], grid[552], grid[553], grid[554], grid[521]);
evolve8 e522 (grid_evolve[522], grid[489], grid[490], grid[491], grid[521], grid[523], grid[553], grid[554], grid[555], grid[522]);
evolve8 e523 (grid_evolve[523], grid[490], grid[491], grid[492], grid[522], grid[524], grid[554], grid[555], grid[556], grid[523]);
evolve8 e524 (grid_evolve[524], grid[491], grid[492], grid[493], grid[523], grid[525], grid[555], grid[556], grid[557], grid[524]);
evolve8 e525 (grid_evolve[525], grid[492], grid[493], grid[494], grid[524], grid[526], grid[556], grid[557], grid[558], grid[525]);
evolve8 e526 (grid_evolve[526], grid[493], grid[494], grid[495], grid[525], grid[527], grid[557], grid[558], grid[559], grid[526]);
evolve8 e527 (grid_evolve[527], grid[494], grid[495], grid[496], grid[526], grid[528], grid[558], grid[559], grid[560], grid[527]);
evolve8 e528 (grid_evolve[528], grid[495], grid[496], grid[497], grid[527], grid[529], grid[559], grid[560], grid[561], grid[528]);
evolve8 e529 (grid_evolve[529], grid[496], grid[497], grid[498], grid[528], grid[530], grid[560], grid[561], grid[562], grid[529]);
evolve8 e530 (grid_evolve[530], grid[497], grid[498], grid[499], grid[529], grid[531], grid[561], grid[562], grid[563], grid[530]);
evolve8 e531 (grid_evolve[531], grid[498], grid[499], grid[500], grid[530], grid[532], grid[562], grid[563], grid[564], grid[531]);
evolve8 e532 (grid_evolve[532], grid[499], grid[500], grid[501], grid[531], grid[533], grid[563], grid[564], grid[565], grid[532]);
evolve8 e533 (grid_evolve[533], grid[500], grid[501], grid[502], grid[532], grid[534], grid[564], grid[565], grid[566], grid[533]);
evolve8 e534 (grid_evolve[534], grid[501], grid[502], grid[503], grid[533], grid[535], grid[565], grid[566], grid[567], grid[534]);
evolve8 e535 (grid_evolve[535], grid[502], grid[503], grid[504], grid[534], grid[536], grid[566], grid[567], grid[568], grid[535]);
evolve8 e536 (grid_evolve[536], grid[503], grid[504], grid[505], grid[535], grid[537], grid[567], grid[568], grid[569], grid[536]);
evolve8 e537 (grid_evolve[537], grid[504], grid[505], grid[506], grid[536], grid[538], grid[568], grid[569], grid[570], grid[537]);
evolve8 e538 (grid_evolve[538], grid[505], grid[506], grid[507], grid[537], grid[539], grid[569], grid[570], grid[571], grid[538]);
evolve8 e539 (grid_evolve[539], grid[506], grid[507], grid[508], grid[538], grid[540], grid[570], grid[571], grid[572], grid[539]);
evolve8 e540 (grid_evolve[540], grid[507], grid[508], grid[509], grid[539], grid[541], grid[571], grid[572], grid[573], grid[540]);
evolve8 e541 (grid_evolve[541], grid[508], grid[509], grid[510], grid[540], grid[542], grid[572], grid[573], grid[574], grid[541]);
evolve8 e542 (grid_evolve[542], grid[509], grid[510], grid[511], grid[541], grid[543], grid[573], grid[574], grid[575], grid[542]);
evolve5 e543 (grid_evolve[543], grid[510], grid[511], grid[542], grid[574], grid[575], grid[543]);

evolve5 e544 (grid_evolve[544], grid[512], grid[513], grid[545], grid[576], grid[577], grid[544]);
evolve8 e545 (grid_evolve[545], grid[512], grid[513], grid[514], grid[544], grid[546], grid[576], grid[577], grid[578], grid[545]);
evolve8 e546 (grid_evolve[546], grid[513], grid[514], grid[515], grid[545], grid[547], grid[577], grid[578], grid[579], grid[546]);
evolve8 e547 (grid_evolve[547], grid[514], grid[515], grid[516], grid[546], grid[548], grid[578], grid[579], grid[580], grid[547]);
evolve8 e548 (grid_evolve[548], grid[515], grid[516], grid[517], grid[547], grid[549], grid[579], grid[580], grid[581], grid[548]);
evolve8 e549 (grid_evolve[549], grid[516], grid[517], grid[518], grid[548], grid[550], grid[580], grid[581], grid[582], grid[549]);
evolve8 e550 (grid_evolve[550], grid[517], grid[518], grid[519], grid[549], grid[551], grid[581], grid[582], grid[583], grid[550]);
evolve8 e551 (grid_evolve[551], grid[518], grid[519], grid[520], grid[550], grid[552], grid[582], grid[583], grid[584], grid[551]);
evolve8 e552 (grid_evolve[552], grid[519], grid[520], grid[521], grid[551], grid[553], grid[583], grid[584], grid[585], grid[552]);
evolve8 e553 (grid_evolve[553], grid[520], grid[521], grid[522], grid[552], grid[554], grid[584], grid[585], grid[586], grid[553]);
evolve8 e554 (grid_evolve[554], grid[521], grid[522], grid[523], grid[553], grid[555], grid[585], grid[586], grid[587], grid[554]);
evolve8 e555 (grid_evolve[555], grid[522], grid[523], grid[524], grid[554], grid[556], grid[586], grid[587], grid[588], grid[555]);
evolve8 e556 (grid_evolve[556], grid[523], grid[524], grid[525], grid[555], grid[557], grid[587], grid[588], grid[589], grid[556]);
evolve8 e557 (grid_evolve[557], grid[524], grid[525], grid[526], grid[556], grid[558], grid[588], grid[589], grid[590], grid[557]);
evolve8 e558 (grid_evolve[558], grid[525], grid[526], grid[527], grid[557], grid[559], grid[589], grid[590], grid[591], grid[558]);
evolve8 e559 (grid_evolve[559], grid[526], grid[527], grid[528], grid[558], grid[560], grid[590], grid[591], grid[592], grid[559]);
evolve8 e560 (grid_evolve[560], grid[527], grid[528], grid[529], grid[559], grid[561], grid[591], grid[592], grid[593], grid[560]);
evolve8 e561 (grid_evolve[561], grid[528], grid[529], grid[530], grid[560], grid[562], grid[592], grid[593], grid[594], grid[561]);
evolve8 e562 (grid_evolve[562], grid[529], grid[530], grid[531], grid[561], grid[563], grid[593], grid[594], grid[595], grid[562]);
evolve8 e563 (grid_evolve[563], grid[530], grid[531], grid[532], grid[562], grid[564], grid[594], grid[595], grid[596], grid[563]);
evolve8 e564 (grid_evolve[564], grid[531], grid[532], grid[533], grid[563], grid[565], grid[595], grid[596], grid[597], grid[564]);
evolve8 e565 (grid_evolve[565], grid[532], grid[533], grid[534], grid[564], grid[566], grid[596], grid[597], grid[598], grid[565]);
evolve8 e566 (grid_evolve[566], grid[533], grid[534], grid[535], grid[565], grid[567], grid[597], grid[598], grid[599], grid[566]);
evolve8 e567 (grid_evolve[567], grid[534], grid[535], grid[536], grid[566], grid[568], grid[598], grid[599], grid[600], grid[567]);
evolve8 e568 (grid_evolve[568], grid[535], grid[536], grid[537], grid[567], grid[569], grid[599], grid[600], grid[601], grid[568]);
evolve8 e569 (grid_evolve[569], grid[536], grid[537], grid[538], grid[568], grid[570], grid[600], grid[601], grid[602], grid[569]);
evolve8 e570 (grid_evolve[570], grid[537], grid[538], grid[539], grid[569], grid[571], grid[601], grid[602], grid[603], grid[570]);
evolve8 e571 (grid_evolve[571], grid[538], grid[539], grid[540], grid[570], grid[572], grid[602], grid[603], grid[604], grid[571]);
evolve8 e572 (grid_evolve[572], grid[539], grid[540], grid[541], grid[571], grid[573], grid[603], grid[604], grid[605], grid[572]);
evolve8 e573 (grid_evolve[573], grid[540], grid[541], grid[542], grid[572], grid[574], grid[604], grid[605], grid[606], grid[573]);
evolve8 e574 (grid_evolve[574], grid[541], grid[542], grid[543], grid[573], grid[575], grid[605], grid[606], grid[607], grid[574]);
evolve5 e575 (grid_evolve[575], grid[542], grid[543], grid[574], grid[606], grid[607], grid[575]);

evolve5 e576 (grid_evolve[576], grid[544], grid[545], grid[577], grid[608], grid[609], grid[576]);
evolve8 e577 (grid_evolve[577], grid[544], grid[545], grid[546], grid[576], grid[578], grid[608], grid[609], grid[610], grid[577]);
evolve8 e578 (grid_evolve[578], grid[545], grid[546], grid[547], grid[577], grid[579], grid[609], grid[610], grid[611], grid[578]);
evolve8 e579 (grid_evolve[579], grid[546], grid[547], grid[548], grid[578], grid[580], grid[610], grid[611], grid[612], grid[579]);
evolve8 e580 (grid_evolve[580], grid[547], grid[548], grid[549], grid[579], grid[581], grid[611], grid[612], grid[613], grid[580]);
evolve8 e581 (grid_evolve[581], grid[548], grid[549], grid[550], grid[580], grid[582], grid[612], grid[613], grid[614], grid[581]);
evolve8 e582 (grid_evolve[582], grid[549], grid[550], grid[551], grid[581], grid[583], grid[613], grid[614], grid[615], grid[582]);
evolve8 e583 (grid_evolve[583], grid[550], grid[551], grid[552], grid[582], grid[584], grid[614], grid[615], grid[616], grid[583]);
evolve8 e584 (grid_evolve[584], grid[551], grid[552], grid[553], grid[583], grid[585], grid[615], grid[616], grid[617], grid[584]);
evolve8 e585 (grid_evolve[585], grid[552], grid[553], grid[554], grid[584], grid[586], grid[616], grid[617], grid[618], grid[585]);
evolve8 e586 (grid_evolve[586], grid[553], grid[554], grid[555], grid[585], grid[587], grid[617], grid[618], grid[619], grid[586]);
evolve8 e587 (grid_evolve[587], grid[554], grid[555], grid[556], grid[586], grid[588], grid[618], grid[619], grid[620], grid[587]);
evolve8 e588 (grid_evolve[588], grid[555], grid[556], grid[557], grid[587], grid[589], grid[619], grid[620], grid[621], grid[588]);
evolve8 e589 (grid_evolve[589], grid[556], grid[557], grid[558], grid[588], grid[590], grid[620], grid[621], grid[622], grid[589]);
evolve8 e590 (grid_evolve[590], grid[557], grid[558], grid[559], grid[589], grid[591], grid[621], grid[622], grid[623], grid[590]);
evolve8 e591 (grid_evolve[591], grid[558], grid[559], grid[560], grid[590], grid[592], grid[622], grid[623], grid[624], grid[591]);
evolve8 e592 (grid_evolve[592], grid[559], grid[560], grid[561], grid[591], grid[593], grid[623], grid[624], grid[625], grid[592]);
evolve8 e593 (grid_evolve[593], grid[560], grid[561], grid[562], grid[592], grid[594], grid[624], grid[625], grid[626], grid[593]);
evolve8 e594 (grid_evolve[594], grid[561], grid[562], grid[563], grid[593], grid[595], grid[625], grid[626], grid[627], grid[594]);
evolve8 e595 (grid_evolve[595], grid[562], grid[563], grid[564], grid[594], grid[596], grid[626], grid[627], grid[628], grid[595]);
evolve8 e596 (grid_evolve[596], grid[563], grid[564], grid[565], grid[595], grid[597], grid[627], grid[628], grid[629], grid[596]);
evolve8 e597 (grid_evolve[597], grid[564], grid[565], grid[566], grid[596], grid[598], grid[628], grid[629], grid[630], grid[597]);
evolve8 e598 (grid_evolve[598], grid[565], grid[566], grid[567], grid[597], grid[599], grid[629], grid[630], grid[631], grid[598]);
evolve8 e599 (grid_evolve[599], grid[566], grid[567], grid[568], grid[598], grid[600], grid[630], grid[631], grid[632], grid[599]);
evolve8 e600 (grid_evolve[600], grid[567], grid[568], grid[569], grid[599], grid[601], grid[631], grid[632], grid[633], grid[600]);
evolve8 e601 (grid_evolve[601], grid[568], grid[569], grid[570], grid[600], grid[602], grid[632], grid[633], grid[634], grid[601]);
evolve8 e602 (grid_evolve[602], grid[569], grid[570], grid[571], grid[601], grid[603], grid[633], grid[634], grid[635], grid[602]);
evolve8 e603 (grid_evolve[603], grid[570], grid[571], grid[572], grid[602], grid[604], grid[634], grid[635], grid[636], grid[603]);
evolve8 e604 (grid_evolve[604], grid[571], grid[572], grid[573], grid[603], grid[605], grid[635], grid[636], grid[637], grid[604]);
evolve8 e605 (grid_evolve[605], grid[572], grid[573], grid[574], grid[604], grid[606], grid[636], grid[637], grid[638], grid[605]);
evolve8 e606 (grid_evolve[606], grid[573], grid[574], grid[575], grid[605], grid[607], grid[637], grid[638], grid[639], grid[606]);
evolve5 e607 (grid_evolve[607], grid[574], grid[575], grid[606], grid[638], grid[639], grid[607]);

evolve5 e608 (grid_evolve[608], grid[576], grid[577], grid[609], grid[640], grid[641], grid[608]);
evolve8 e609 (grid_evolve[609], grid[576], grid[577], grid[578], grid[608], grid[610], grid[640], grid[641], grid[642], grid[609]);
evolve8 e610 (grid_evolve[610], grid[577], grid[578], grid[579], grid[609], grid[611], grid[641], grid[642], grid[643], grid[610]);
evolve8 e611 (grid_evolve[611], grid[578], grid[579], grid[580], grid[610], grid[612], grid[642], grid[643], grid[644], grid[611]);
evolve8 e612 (grid_evolve[612], grid[579], grid[580], grid[581], grid[611], grid[613], grid[643], grid[644], grid[645], grid[612]);
evolve8 e613 (grid_evolve[613], grid[580], grid[581], grid[582], grid[612], grid[614], grid[644], grid[645], grid[646], grid[613]);
evolve8 e614 (grid_evolve[614], grid[581], grid[582], grid[583], grid[613], grid[615], grid[645], grid[646], grid[647], grid[614]);
evolve8 e615 (grid_evolve[615], grid[582], grid[583], grid[584], grid[614], grid[616], grid[646], grid[647], grid[648], grid[615]);
evolve8 e616 (grid_evolve[616], grid[583], grid[584], grid[585], grid[615], grid[617], grid[647], grid[648], grid[649], grid[616]);
evolve8 e617 (grid_evolve[617], grid[584], grid[585], grid[586], grid[616], grid[618], grid[648], grid[649], grid[650], grid[617]);
evolve8 e618 (grid_evolve[618], grid[585], grid[586], grid[587], grid[617], grid[619], grid[649], grid[650], grid[651], grid[618]);
evolve8 e619 (grid_evolve[619], grid[586], grid[587], grid[588], grid[618], grid[620], grid[650], grid[651], grid[652], grid[619]);
evolve8 e620 (grid_evolve[620], grid[587], grid[588], grid[589], grid[619], grid[621], grid[651], grid[652], grid[653], grid[620]);
evolve8 e621 (grid_evolve[621], grid[588], grid[589], grid[590], grid[620], grid[622], grid[652], grid[653], grid[654], grid[621]);
evolve8 e622 (grid_evolve[622], grid[589], grid[590], grid[591], grid[621], grid[623], grid[653], grid[654], grid[655], grid[622]);
evolve8 e623 (grid_evolve[623], grid[590], grid[591], grid[592], grid[622], grid[624], grid[654], grid[655], grid[656], grid[623]);
evolve8 e624 (grid_evolve[624], grid[591], grid[592], grid[593], grid[623], grid[625], grid[655], grid[656], grid[657], grid[624]);
evolve8 e625 (grid_evolve[625], grid[592], grid[593], grid[594], grid[624], grid[626], grid[656], grid[657], grid[658], grid[625]);
evolve8 e626 (grid_evolve[626], grid[593], grid[594], grid[595], grid[625], grid[627], grid[657], grid[658], grid[659], grid[626]);
evolve8 e627 (grid_evolve[627], grid[594], grid[595], grid[596], grid[626], grid[628], grid[658], grid[659], grid[660], grid[627]);
evolve8 e628 (grid_evolve[628], grid[595], grid[596], grid[597], grid[627], grid[629], grid[659], grid[660], grid[661], grid[628]);
evolve8 e629 (grid_evolve[629], grid[596], grid[597], grid[598], grid[628], grid[630], grid[660], grid[661], grid[662], grid[629]);
evolve8 e630 (grid_evolve[630], grid[597], grid[598], grid[599], grid[629], grid[631], grid[661], grid[662], grid[663], grid[630]);
evolve8 e631 (grid_evolve[631], grid[598], grid[599], grid[600], grid[630], grid[632], grid[662], grid[663], grid[664], grid[631]);
evolve8 e632 (grid_evolve[632], grid[599], grid[600], grid[601], grid[631], grid[633], grid[663], grid[664], grid[665], grid[632]);
evolve8 e633 (grid_evolve[633], grid[600], grid[601], grid[602], grid[632], grid[634], grid[664], grid[665], grid[666], grid[633]);
evolve8 e634 (grid_evolve[634], grid[601], grid[602], grid[603], grid[633], grid[635], grid[665], grid[666], grid[667], grid[634]);
evolve8 e635 (grid_evolve[635], grid[602], grid[603], grid[604], grid[634], grid[636], grid[666], grid[667], grid[668], grid[635]);
evolve8 e636 (grid_evolve[636], grid[603], grid[604], grid[605], grid[635], grid[637], grid[667], grid[668], grid[669], grid[636]);
evolve8 e637 (grid_evolve[637], grid[604], grid[605], grid[606], grid[636], grid[638], grid[668], grid[669], grid[670], grid[637]);
evolve8 e638 (grid_evolve[638], grid[605], grid[606], grid[607], grid[637], grid[639], grid[669], grid[670], grid[671], grid[638]);
evolve5 e639 (grid_evolve[639], grid[606], grid[607], grid[638], grid[670], grid[671], grid[639]);

evolve5 e640 (grid_evolve[640], grid[608], grid[609], grid[641], grid[672], grid[673], grid[640]);
evolve8 e641 (grid_evolve[641], grid[608], grid[609], grid[610], grid[640], grid[642], grid[672], grid[673], grid[674], grid[641]);
evolve8 e642 (grid_evolve[642], grid[609], grid[610], grid[611], grid[641], grid[643], grid[673], grid[674], grid[675], grid[642]);
evolve8 e643 (grid_evolve[643], grid[610], grid[611], grid[612], grid[642], grid[644], grid[674], grid[675], grid[676], grid[643]);
evolve8 e644 (grid_evolve[644], grid[611], grid[612], grid[613], grid[643], grid[645], grid[675], grid[676], grid[677], grid[644]);
evolve8 e645 (grid_evolve[645], grid[612], grid[613], grid[614], grid[644], grid[646], grid[676], grid[677], grid[678], grid[645]);
evolve8 e646 (grid_evolve[646], grid[613], grid[614], grid[615], grid[645], grid[647], grid[677], grid[678], grid[679], grid[646]);
evolve8 e647 (grid_evolve[647], grid[614], grid[615], grid[616], grid[646], grid[648], grid[678], grid[679], grid[680], grid[647]);
evolve8 e648 (grid_evolve[648], grid[615], grid[616], grid[617], grid[647], grid[649], grid[679], grid[680], grid[681], grid[648]);
evolve8 e649 (grid_evolve[649], grid[616], grid[617], grid[618], grid[648], grid[650], grid[680], grid[681], grid[682], grid[649]);
evolve8 e650 (grid_evolve[650], grid[617], grid[618], grid[619], grid[649], grid[651], grid[681], grid[682], grid[683], grid[650]);
evolve8 e651 (grid_evolve[651], grid[618], grid[619], grid[620], grid[650], grid[652], grid[682], grid[683], grid[684], grid[651]);
evolve8 e652 (grid_evolve[652], grid[619], grid[620], grid[621], grid[651], grid[653], grid[683], grid[684], grid[685], grid[652]);
evolve8 e653 (grid_evolve[653], grid[620], grid[621], grid[622], grid[652], grid[654], grid[684], grid[685], grid[686], grid[653]);
evolve8 e654 (grid_evolve[654], grid[621], grid[622], grid[623], grid[653], grid[655], grid[685], grid[686], grid[687], grid[654]);
evolve8 e655 (grid_evolve[655], grid[622], grid[623], grid[624], grid[654], grid[656], grid[686], grid[687], grid[688], grid[655]);
evolve8 e656 (grid_evolve[656], grid[623], grid[624], grid[625], grid[655], grid[657], grid[687], grid[688], grid[689], grid[656]);
evolve8 e657 (grid_evolve[657], grid[624], grid[625], grid[626], grid[656], grid[658], grid[688], grid[689], grid[690], grid[657]);
evolve8 e658 (grid_evolve[658], grid[625], grid[626], grid[627], grid[657], grid[659], grid[689], grid[690], grid[691], grid[658]);
evolve8 e659 (grid_evolve[659], grid[626], grid[627], grid[628], grid[658], grid[660], grid[690], grid[691], grid[692], grid[659]);
evolve8 e660 (grid_evolve[660], grid[627], grid[628], grid[629], grid[659], grid[661], grid[691], grid[692], grid[693], grid[660]);
evolve8 e661 (grid_evolve[661], grid[628], grid[629], grid[630], grid[660], grid[662], grid[692], grid[693], grid[694], grid[661]);
evolve8 e662 (grid_evolve[662], grid[629], grid[630], grid[631], grid[661], grid[663], grid[693], grid[694], grid[695], grid[662]);
evolve8 e663 (grid_evolve[663], grid[630], grid[631], grid[632], grid[662], grid[664], grid[694], grid[695], grid[696], grid[663]);
evolve8 e664 (grid_evolve[664], grid[631], grid[632], grid[633], grid[663], grid[665], grid[695], grid[696], grid[697], grid[664]);
evolve8 e665 (grid_evolve[665], grid[632], grid[633], grid[634], grid[664], grid[666], grid[696], grid[697], grid[698], grid[665]);
evolve8 e666 (grid_evolve[666], grid[633], grid[634], grid[635], grid[665], grid[667], grid[697], grid[698], grid[699], grid[666]);
evolve8 e667 (grid_evolve[667], grid[634], grid[635], grid[636], grid[666], grid[668], grid[698], grid[699], grid[700], grid[667]);
evolve8 e668 (grid_evolve[668], grid[635], grid[636], grid[637], grid[667], grid[669], grid[699], grid[700], grid[701], grid[668]);
evolve8 e669 (grid_evolve[669], grid[636], grid[637], grid[638], grid[668], grid[670], grid[700], grid[701], grid[702], grid[669]);
evolve8 e670 (grid_evolve[670], grid[637], grid[638], grid[639], grid[669], grid[671], grid[701], grid[702], grid[703], grid[670]);
evolve5 e671 (grid_evolve[671], grid[638], grid[639], grid[670], grid[702], grid[703], grid[671]);

evolve5 e672 (grid_evolve[672], grid[640], grid[641], grid[673], grid[704], grid[705], grid[672]);
evolve8 e673 (grid_evolve[673], grid[640], grid[641], grid[642], grid[672], grid[674], grid[704], grid[705], grid[706], grid[673]);
evolve8 e674 (grid_evolve[674], grid[641], grid[642], grid[643], grid[673], grid[675], grid[705], grid[706], grid[707], grid[674]);
evolve8 e675 (grid_evolve[675], grid[642], grid[643], grid[644], grid[674], grid[676], grid[706], grid[707], grid[708], grid[675]);
evolve8 e676 (grid_evolve[676], grid[643], grid[644], grid[645], grid[675], grid[677], grid[707], grid[708], grid[709], grid[676]);
evolve8 e677 (grid_evolve[677], grid[644], grid[645], grid[646], grid[676], grid[678], grid[708], grid[709], grid[710], grid[677]);
evolve8 e678 (grid_evolve[678], grid[645], grid[646], grid[647], grid[677], grid[679], grid[709], grid[710], grid[711], grid[678]);
evolve8 e679 (grid_evolve[679], grid[646], grid[647], grid[648], grid[678], grid[680], grid[710], grid[711], grid[712], grid[679]);
evolve8 e680 (grid_evolve[680], grid[647], grid[648], grid[649], grid[679], grid[681], grid[711], grid[712], grid[713], grid[680]);
evolve8 e681 (grid_evolve[681], grid[648], grid[649], grid[650], grid[680], grid[682], grid[712], grid[713], grid[714], grid[681]);
evolve8 e682 (grid_evolve[682], grid[649], grid[650], grid[651], grid[681], grid[683], grid[713], grid[714], grid[715], grid[682]);
evolve8 e683 (grid_evolve[683], grid[650], grid[651], grid[652], grid[682], grid[684], grid[714], grid[715], grid[716], grid[683]);
evolve8 e684 (grid_evolve[684], grid[651], grid[652], grid[653], grid[683], grid[685], grid[715], grid[716], grid[717], grid[684]);
evolve8 e685 (grid_evolve[685], grid[652], grid[653], grid[654], grid[684], grid[686], grid[716], grid[717], grid[718], grid[685]);
evolve8 e686 (grid_evolve[686], grid[653], grid[654], grid[655], grid[685], grid[687], grid[717], grid[718], grid[719], grid[686]);
evolve8 e687 (grid_evolve[687], grid[654], grid[655], grid[656], grid[686], grid[688], grid[718], grid[719], grid[720], grid[687]);
evolve8 e688 (grid_evolve[688], grid[655], grid[656], grid[657], grid[687], grid[689], grid[719], grid[720], grid[721], grid[688]);
evolve8 e689 (grid_evolve[689], grid[656], grid[657], grid[658], grid[688], grid[690], grid[720], grid[721], grid[722], grid[689]);
evolve8 e690 (grid_evolve[690], grid[657], grid[658], grid[659], grid[689], grid[691], grid[721], grid[722], grid[723], grid[690]);
evolve8 e691 (grid_evolve[691], grid[658], grid[659], grid[660], grid[690], grid[692], grid[722], grid[723], grid[724], grid[691]);
evolve8 e692 (grid_evolve[692], grid[659], grid[660], grid[661], grid[691], grid[693], grid[723], grid[724], grid[725], grid[692]);
evolve8 e693 (grid_evolve[693], grid[660], grid[661], grid[662], grid[692], grid[694], grid[724], grid[725], grid[726], grid[693]);
evolve8 e694 (grid_evolve[694], grid[661], grid[662], grid[663], grid[693], grid[695], grid[725], grid[726], grid[727], grid[694]);
evolve8 e695 (grid_evolve[695], grid[662], grid[663], grid[664], grid[694], grid[696], grid[726], grid[727], grid[728], grid[695]);
evolve8 e696 (grid_evolve[696], grid[663], grid[664], grid[665], grid[695], grid[697], grid[727], grid[728], grid[729], grid[696]);
evolve8 e697 (grid_evolve[697], grid[664], grid[665], grid[666], grid[696], grid[698], grid[728], grid[729], grid[730], grid[697]);
evolve8 e698 (grid_evolve[698], grid[665], grid[666], grid[667], grid[697], grid[699], grid[729], grid[730], grid[731], grid[698]);
evolve8 e699 (grid_evolve[699], grid[666], grid[667], grid[668], grid[698], grid[700], grid[730], grid[731], grid[732], grid[699]);
evolve8 e700 (grid_evolve[700], grid[667], grid[668], grid[669], grid[699], grid[701], grid[731], grid[732], grid[733], grid[700]);
evolve8 e701 (grid_evolve[701], grid[668], grid[669], grid[670], grid[700], grid[702], grid[732], grid[733], grid[734], grid[701]);
evolve8 e702 (grid_evolve[702], grid[669], grid[670], grid[671], grid[701], grid[703], grid[733], grid[734], grid[735], grid[702]);
evolve5 e703 (grid_evolve[703], grid[670], grid[671], grid[702], grid[734], grid[735], grid[703]);

evolve5 e704 (grid_evolve[704], grid[672], grid[673], grid[705], grid[736], grid[737], grid[704]);
evolve8 e705 (grid_evolve[705], grid[672], grid[673], grid[674], grid[704], grid[706], grid[736], grid[737], grid[738], grid[705]);
evolve8 e706 (grid_evolve[706], grid[673], grid[674], grid[675], grid[705], grid[707], grid[737], grid[738], grid[739], grid[706]);
evolve8 e707 (grid_evolve[707], grid[674], grid[675], grid[676], grid[706], grid[708], grid[738], grid[739], grid[740], grid[707]);
evolve8 e708 (grid_evolve[708], grid[675], grid[676], grid[677], grid[707], grid[709], grid[739], grid[740], grid[741], grid[708]);
evolve8 e709 (grid_evolve[709], grid[676], grid[677], grid[678], grid[708], grid[710], grid[740], grid[741], grid[742], grid[709]);
evolve8 e710 (grid_evolve[710], grid[677], grid[678], grid[679], grid[709], grid[711], grid[741], grid[742], grid[743], grid[710]);
evolve8 e711 (grid_evolve[711], grid[678], grid[679], grid[680], grid[710], grid[712], grid[742], grid[743], grid[744], grid[711]);
evolve8 e712 (grid_evolve[712], grid[679], grid[680], grid[681], grid[711], grid[713], grid[743], grid[744], grid[745], grid[712]);
evolve8 e713 (grid_evolve[713], grid[680], grid[681], grid[682], grid[712], grid[714], grid[744], grid[745], grid[746], grid[713]);
evolve8 e714 (grid_evolve[714], grid[681], grid[682], grid[683], grid[713], grid[715], grid[745], grid[746], grid[747], grid[714]);
evolve8 e715 (grid_evolve[715], grid[682], grid[683], grid[684], grid[714], grid[716], grid[746], grid[747], grid[748], grid[715]);
evolve8 e716 (grid_evolve[716], grid[683], grid[684], grid[685], grid[715], grid[717], grid[747], grid[748], grid[749], grid[716]);
evolve8 e717 (grid_evolve[717], grid[684], grid[685], grid[686], grid[716], grid[718], grid[748], grid[749], grid[750], grid[717]);
evolve8 e718 (grid_evolve[718], grid[685], grid[686], grid[687], grid[717], grid[719], grid[749], grid[750], grid[751], grid[718]);
evolve8 e719 (grid_evolve[719], grid[686], grid[687], grid[688], grid[718], grid[720], grid[750], grid[751], grid[752], grid[719]);
evolve8 e720 (grid_evolve[720], grid[687], grid[688], grid[689], grid[719], grid[721], grid[751], grid[752], grid[753], grid[720]);
evolve8 e721 (grid_evolve[721], grid[688], grid[689], grid[690], grid[720], grid[722], grid[752], grid[753], grid[754], grid[721]);
evolve8 e722 (grid_evolve[722], grid[689], grid[690], grid[691], grid[721], grid[723], grid[753], grid[754], grid[755], grid[722]);
evolve8 e723 (grid_evolve[723], grid[690], grid[691], grid[692], grid[722], grid[724], grid[754], grid[755], grid[756], grid[723]);
evolve8 e724 (grid_evolve[724], grid[691], grid[692], grid[693], grid[723], grid[725], grid[755], grid[756], grid[757], grid[724]);
evolve8 e725 (grid_evolve[725], grid[692], grid[693], grid[694], grid[724], grid[726], grid[756], grid[757], grid[758], grid[725]);
evolve8 e726 (grid_evolve[726], grid[693], grid[694], grid[695], grid[725], grid[727], grid[757], grid[758], grid[759], grid[726]);
evolve8 e727 (grid_evolve[727], grid[694], grid[695], grid[696], grid[726], grid[728], grid[758], grid[759], grid[760], grid[727]);
evolve8 e728 (grid_evolve[728], grid[695], grid[696], grid[697], grid[727], grid[729], grid[759], grid[760], grid[761], grid[728]);
evolve8 e729 (grid_evolve[729], grid[696], grid[697], grid[698], grid[728], grid[730], grid[760], grid[761], grid[762], grid[729]);
evolve8 e730 (grid_evolve[730], grid[697], grid[698], grid[699], grid[729], grid[731], grid[761], grid[762], grid[763], grid[730]);
evolve8 e731 (grid_evolve[731], grid[698], grid[699], grid[700], grid[730], grid[732], grid[762], grid[763], grid[764], grid[731]);
evolve8 e732 (grid_evolve[732], grid[699], grid[700], grid[701], grid[731], grid[733], grid[763], grid[764], grid[765], grid[732]);
evolve8 e733 (grid_evolve[733], grid[700], grid[701], grid[702], grid[732], grid[734], grid[764], grid[765], grid[766], grid[733]);
evolve8 e734 (grid_evolve[734], grid[701], grid[702], grid[703], grid[733], grid[735], grid[765], grid[766], grid[767], grid[734]);
evolve5 e735 (grid_evolve[735], grid[702], grid[703], grid[734], grid[766], grid[767], grid[735]);

evolve5 e736 (grid_evolve[736], grid[704], grid[705], grid[737], grid[768], grid[769], grid[736]);
evolve8 e737 (grid_evolve[737], grid[704], grid[705], grid[706], grid[736], grid[738], grid[768], grid[769], grid[770], grid[737]);
evolve8 e738 (grid_evolve[738], grid[705], grid[706], grid[707], grid[737], grid[739], grid[769], grid[770], grid[771], grid[738]);
evolve8 e739 (grid_evolve[739], grid[706], grid[707], grid[708], grid[738], grid[740], grid[770], grid[771], grid[772], grid[739]);
evolve8 e740 (grid_evolve[740], grid[707], grid[708], grid[709], grid[739], grid[741], grid[771], grid[772], grid[773], grid[740]);
evolve8 e741 (grid_evolve[741], grid[708], grid[709], grid[710], grid[740], grid[742], grid[772], grid[773], grid[774], grid[741]);
evolve8 e742 (grid_evolve[742], grid[709], grid[710], grid[711], grid[741], grid[743], grid[773], grid[774], grid[775], grid[742]);
evolve8 e743 (grid_evolve[743], grid[710], grid[711], grid[712], grid[742], grid[744], grid[774], grid[775], grid[776], grid[743]);
evolve8 e744 (grid_evolve[744], grid[711], grid[712], grid[713], grid[743], grid[745], grid[775], grid[776], grid[777], grid[744]);
evolve8 e745 (grid_evolve[745], grid[712], grid[713], grid[714], grid[744], grid[746], grid[776], grid[777], grid[778], grid[745]);
evolve8 e746 (grid_evolve[746], grid[713], grid[714], grid[715], grid[745], grid[747], grid[777], grid[778], grid[779], grid[746]);
evolve8 e747 (grid_evolve[747], grid[714], grid[715], grid[716], grid[746], grid[748], grid[778], grid[779], grid[780], grid[747]);
evolve8 e748 (grid_evolve[748], grid[715], grid[716], grid[717], grid[747], grid[749], grid[779], grid[780], grid[781], grid[748]);
evolve8 e749 (grid_evolve[749], grid[716], grid[717], grid[718], grid[748], grid[750], grid[780], grid[781], grid[782], grid[749]);
evolve8 e750 (grid_evolve[750], grid[717], grid[718], grid[719], grid[749], grid[751], grid[781], grid[782], grid[783], grid[750]);
evolve8 e751 (grid_evolve[751], grid[718], grid[719], grid[720], grid[750], grid[752], grid[782], grid[783], grid[784], grid[751]);
evolve8 e752 (grid_evolve[752], grid[719], grid[720], grid[721], grid[751], grid[753], grid[783], grid[784], grid[785], grid[752]);
evolve8 e753 (grid_evolve[753], grid[720], grid[721], grid[722], grid[752], grid[754], grid[784], grid[785], grid[786], grid[753]);
evolve8 e754 (grid_evolve[754], grid[721], grid[722], grid[723], grid[753], grid[755], grid[785], grid[786], grid[787], grid[754]);
evolve8 e755 (grid_evolve[755], grid[722], grid[723], grid[724], grid[754], grid[756], grid[786], grid[787], grid[788], grid[755]);
evolve8 e756 (grid_evolve[756], grid[723], grid[724], grid[725], grid[755], grid[757], grid[787], grid[788], grid[789], grid[756]);
evolve8 e757 (grid_evolve[757], grid[724], grid[725], grid[726], grid[756], grid[758], grid[788], grid[789], grid[790], grid[757]);
evolve8 e758 (grid_evolve[758], grid[725], grid[726], grid[727], grid[757], grid[759], grid[789], grid[790], grid[791], grid[758]);
evolve8 e759 (grid_evolve[759], grid[726], grid[727], grid[728], grid[758], grid[760], grid[790], grid[791], grid[792], grid[759]);
evolve8 e760 (grid_evolve[760], grid[727], grid[728], grid[729], grid[759], grid[761], grid[791], grid[792], grid[793], grid[760]);
evolve8 e761 (grid_evolve[761], grid[728], grid[729], grid[730], grid[760], grid[762], grid[792], grid[793], grid[794], grid[761]);
evolve8 e762 (grid_evolve[762], grid[729], grid[730], grid[731], grid[761], grid[763], grid[793], grid[794], grid[795], grid[762]);
evolve8 e763 (grid_evolve[763], grid[730], grid[731], grid[732], grid[762], grid[764], grid[794], grid[795], grid[796], grid[763]);
evolve8 e764 (grid_evolve[764], grid[731], grid[732], grid[733], grid[763], grid[765], grid[795], grid[796], grid[797], grid[764]);
evolve8 e765 (grid_evolve[765], grid[732], grid[733], grid[734], grid[764], grid[766], grid[796], grid[797], grid[798], grid[765]);
evolve8 e766 (grid_evolve[766], grid[733], grid[734], grid[735], grid[765], grid[767], grid[797], grid[798], grid[799], grid[766]);
evolve5 e767 (grid_evolve[767], grid[734], grid[735], grid[766], grid[798], grid[799], grid[767]);

evolve5 e768 (grid_evolve[768], grid[736], grid[737], grid[769], grid[800], grid[801], grid[768]);
evolve8 e769 (grid_evolve[769], grid[736], grid[737], grid[738], grid[768], grid[770], grid[800], grid[801], grid[802], grid[769]);
evolve8 e770 (grid_evolve[770], grid[737], grid[738], grid[739], grid[769], grid[771], grid[801], grid[802], grid[803], grid[770]);
evolve8 e771 (grid_evolve[771], grid[738], grid[739], grid[740], grid[770], grid[772], grid[802], grid[803], grid[804], grid[771]);
evolve8 e772 (grid_evolve[772], grid[739], grid[740], grid[741], grid[771], grid[773], grid[803], grid[804], grid[805], grid[772]);
evolve8 e773 (grid_evolve[773], grid[740], grid[741], grid[742], grid[772], grid[774], grid[804], grid[805], grid[806], grid[773]);
evolve8 e774 (grid_evolve[774], grid[741], grid[742], grid[743], grid[773], grid[775], grid[805], grid[806], grid[807], grid[774]);
evolve8 e775 (grid_evolve[775], grid[742], grid[743], grid[744], grid[774], grid[776], grid[806], grid[807], grid[808], grid[775]);
evolve8 e776 (grid_evolve[776], grid[743], grid[744], grid[745], grid[775], grid[777], grid[807], grid[808], grid[809], grid[776]);
evolve8 e777 (grid_evolve[777], grid[744], grid[745], grid[746], grid[776], grid[778], grid[808], grid[809], grid[810], grid[777]);
evolve8 e778 (grid_evolve[778], grid[745], grid[746], grid[747], grid[777], grid[779], grid[809], grid[810], grid[811], grid[778]);
evolve8 e779 (grid_evolve[779], grid[746], grid[747], grid[748], grid[778], grid[780], grid[810], grid[811], grid[812], grid[779]);
evolve8 e780 (grid_evolve[780], grid[747], grid[748], grid[749], grid[779], grid[781], grid[811], grid[812], grid[813], grid[780]);
evolve8 e781 (grid_evolve[781], grid[748], grid[749], grid[750], grid[780], grid[782], grid[812], grid[813], grid[814], grid[781]);
evolve8 e782 (grid_evolve[782], grid[749], grid[750], grid[751], grid[781], grid[783], grid[813], grid[814], grid[815], grid[782]);
evolve8 e783 (grid_evolve[783], grid[750], grid[751], grid[752], grid[782], grid[784], grid[814], grid[815], grid[816], grid[783]);
evolve8 e784 (grid_evolve[784], grid[751], grid[752], grid[753], grid[783], grid[785], grid[815], grid[816], grid[817], grid[784]);
evolve8 e785 (grid_evolve[785], grid[752], grid[753], grid[754], grid[784], grid[786], grid[816], grid[817], grid[818], grid[785]);
evolve8 e786 (grid_evolve[786], grid[753], grid[754], grid[755], grid[785], grid[787], grid[817], grid[818], grid[819], grid[786]);
evolve8 e787 (grid_evolve[787], grid[754], grid[755], grid[756], grid[786], grid[788], grid[818], grid[819], grid[820], grid[787]);
evolve8 e788 (grid_evolve[788], grid[755], grid[756], grid[757], grid[787], grid[789], grid[819], grid[820], grid[821], grid[788]);
evolve8 e789 (grid_evolve[789], grid[756], grid[757], grid[758], grid[788], grid[790], grid[820], grid[821], grid[822], grid[789]);
evolve8 e790 (grid_evolve[790], grid[757], grid[758], grid[759], grid[789], grid[791], grid[821], grid[822], grid[823], grid[790]);
evolve8 e791 (grid_evolve[791], grid[758], grid[759], grid[760], grid[790], grid[792], grid[822], grid[823], grid[824], grid[791]);
evolve8 e792 (grid_evolve[792], grid[759], grid[760], grid[761], grid[791], grid[793], grid[823], grid[824], grid[825], grid[792]);
evolve8 e793 (grid_evolve[793], grid[760], grid[761], grid[762], grid[792], grid[794], grid[824], grid[825], grid[826], grid[793]);
evolve8 e794 (grid_evolve[794], grid[761], grid[762], grid[763], grid[793], grid[795], grid[825], grid[826], grid[827], grid[794]);
evolve8 e795 (grid_evolve[795], grid[762], grid[763], grid[764], grid[794], grid[796], grid[826], grid[827], grid[828], grid[795]);
evolve8 e796 (grid_evolve[796], grid[763], grid[764], grid[765], grid[795], grid[797], grid[827], grid[828], grid[829], grid[796]);
evolve8 e797 (grid_evolve[797], grid[764], grid[765], grid[766], grid[796], grid[798], grid[828], grid[829], grid[830], grid[797]);
evolve8 e798 (grid_evolve[798], grid[765], grid[766], grid[767], grid[797], grid[799], grid[829], grid[830], grid[831], grid[798]);
evolve5 e799 (grid_evolve[799], grid[766], grid[767], grid[798], grid[830], grid[831], grid[799]);

evolve5 e800 (grid_evolve[800], grid[768], grid[769], grid[801], grid[832], grid[833], grid[800]);
evolve8 e801 (grid_evolve[801], grid[768], grid[769], grid[770], grid[800], grid[802], grid[832], grid[833], grid[834], grid[801]);
evolve8 e802 (grid_evolve[802], grid[769], grid[770], grid[771], grid[801], grid[803], grid[833], grid[834], grid[835], grid[802]);
evolve8 e803 (grid_evolve[803], grid[770], grid[771], grid[772], grid[802], grid[804], grid[834], grid[835], grid[836], grid[803]);
evolve8 e804 (grid_evolve[804], grid[771], grid[772], grid[773], grid[803], grid[805], grid[835], grid[836], grid[837], grid[804]);
evolve8 e805 (grid_evolve[805], grid[772], grid[773], grid[774], grid[804], grid[806], grid[836], grid[837], grid[838], grid[805]);
evolve8 e806 (grid_evolve[806], grid[773], grid[774], grid[775], grid[805], grid[807], grid[837], grid[838], grid[839], grid[806]);
evolve8 e807 (grid_evolve[807], grid[774], grid[775], grid[776], grid[806], grid[808], grid[838], grid[839], grid[840], grid[807]);
evolve8 e808 (grid_evolve[808], grid[775], grid[776], grid[777], grid[807], grid[809], grid[839], grid[840], grid[841], grid[808]);
evolve8 e809 (grid_evolve[809], grid[776], grid[777], grid[778], grid[808], grid[810], grid[840], grid[841], grid[842], grid[809]);
evolve8 e810 (grid_evolve[810], grid[777], grid[778], grid[779], grid[809], grid[811], grid[841], grid[842], grid[843], grid[810]);
evolve8 e811 (grid_evolve[811], grid[778], grid[779], grid[780], grid[810], grid[812], grid[842], grid[843], grid[844], grid[811]);
evolve8 e812 (grid_evolve[812], grid[779], grid[780], grid[781], grid[811], grid[813], grid[843], grid[844], grid[845], grid[812]);
evolve8 e813 (grid_evolve[813], grid[780], grid[781], grid[782], grid[812], grid[814], grid[844], grid[845], grid[846], grid[813]);
evolve8 e814 (grid_evolve[814], grid[781], grid[782], grid[783], grid[813], grid[815], grid[845], grid[846], grid[847], grid[814]);
evolve8 e815 (grid_evolve[815], grid[782], grid[783], grid[784], grid[814], grid[816], grid[846], grid[847], grid[848], grid[815]);
evolve8 e816 (grid_evolve[816], grid[783], grid[784], grid[785], grid[815], grid[817], grid[847], grid[848], grid[849], grid[816]);
evolve8 e817 (grid_evolve[817], grid[784], grid[785], grid[786], grid[816], grid[818], grid[848], grid[849], grid[850], grid[817]);
evolve8 e818 (grid_evolve[818], grid[785], grid[786], grid[787], grid[817], grid[819], grid[849], grid[850], grid[851], grid[818]);
evolve8 e819 (grid_evolve[819], grid[786], grid[787], grid[788], grid[818], grid[820], grid[850], grid[851], grid[852], grid[819]);
evolve8 e820 (grid_evolve[820], grid[787], grid[788], grid[789], grid[819], grid[821], grid[851], grid[852], grid[853], grid[820]);
evolve8 e821 (grid_evolve[821], grid[788], grid[789], grid[790], grid[820], grid[822], grid[852], grid[853], grid[854], grid[821]);
evolve8 e822 (grid_evolve[822], grid[789], grid[790], grid[791], grid[821], grid[823], grid[853], grid[854], grid[855], grid[822]);
evolve8 e823 (grid_evolve[823], grid[790], grid[791], grid[792], grid[822], grid[824], grid[854], grid[855], grid[856], grid[823]);
evolve8 e824 (grid_evolve[824], grid[791], grid[792], grid[793], grid[823], grid[825], grid[855], grid[856], grid[857], grid[824]);
evolve8 e825 (grid_evolve[825], grid[792], grid[793], grid[794], grid[824], grid[826], grid[856], grid[857], grid[858], grid[825]);
evolve8 e826 (grid_evolve[826], grid[793], grid[794], grid[795], grid[825], grid[827], grid[857], grid[858], grid[859], grid[826]);
evolve8 e827 (grid_evolve[827], grid[794], grid[795], grid[796], grid[826], grid[828], grid[858], grid[859], grid[860], grid[827]);
evolve8 e828 (grid_evolve[828], grid[795], grid[796], grid[797], grid[827], grid[829], grid[859], grid[860], grid[861], grid[828]);
evolve8 e829 (grid_evolve[829], grid[796], grid[797], grid[798], grid[828], grid[830], grid[860], grid[861], grid[862], grid[829]);
evolve8 e830 (grid_evolve[830], grid[797], grid[798], grid[799], grid[829], grid[831], grid[861], grid[862], grid[863], grid[830]);
evolve5 e831 (grid_evolve[831], grid[798], grid[799], grid[830], grid[862], grid[863], grid[831]);

evolve5 e832 (grid_evolve[832], grid[800], grid[801], grid[833], grid[864], grid[865], grid[832]);
evolve8 e833 (grid_evolve[833], grid[800], grid[801], grid[802], grid[832], grid[834], grid[864], grid[865], grid[866], grid[833]);
evolve8 e834 (grid_evolve[834], grid[801], grid[802], grid[803], grid[833], grid[835], grid[865], grid[866], grid[867], grid[834]);
evolve8 e835 (grid_evolve[835], grid[802], grid[803], grid[804], grid[834], grid[836], grid[866], grid[867], grid[868], grid[835]);
evolve8 e836 (grid_evolve[836], grid[803], grid[804], grid[805], grid[835], grid[837], grid[867], grid[868], grid[869], grid[836]);
evolve8 e837 (grid_evolve[837], grid[804], grid[805], grid[806], grid[836], grid[838], grid[868], grid[869], grid[870], grid[837]);
evolve8 e838 (grid_evolve[838], grid[805], grid[806], grid[807], grid[837], grid[839], grid[869], grid[870], grid[871], grid[838]);
evolve8 e839 (grid_evolve[839], grid[806], grid[807], grid[808], grid[838], grid[840], grid[870], grid[871], grid[872], grid[839]);
evolve8 e840 (grid_evolve[840], grid[807], grid[808], grid[809], grid[839], grid[841], grid[871], grid[872], grid[873], grid[840]);
evolve8 e841 (grid_evolve[841], grid[808], grid[809], grid[810], grid[840], grid[842], grid[872], grid[873], grid[874], grid[841]);
evolve8 e842 (grid_evolve[842], grid[809], grid[810], grid[811], grid[841], grid[843], grid[873], grid[874], grid[875], grid[842]);
evolve8 e843 (grid_evolve[843], grid[810], grid[811], grid[812], grid[842], grid[844], grid[874], grid[875], grid[876], grid[843]);
evolve8 e844 (grid_evolve[844], grid[811], grid[812], grid[813], grid[843], grid[845], grid[875], grid[876], grid[877], grid[844]);
evolve8 e845 (grid_evolve[845], grid[812], grid[813], grid[814], grid[844], grid[846], grid[876], grid[877], grid[878], grid[845]);
evolve8 e846 (grid_evolve[846], grid[813], grid[814], grid[815], grid[845], grid[847], grid[877], grid[878], grid[879], grid[846]);
evolve8 e847 (grid_evolve[847], grid[814], grid[815], grid[816], grid[846], grid[848], grid[878], grid[879], grid[880], grid[847]);
evolve8 e848 (grid_evolve[848], grid[815], grid[816], grid[817], grid[847], grid[849], grid[879], grid[880], grid[881], grid[848]);
evolve8 e849 (grid_evolve[849], grid[816], grid[817], grid[818], grid[848], grid[850], grid[880], grid[881], grid[882], grid[849]);
evolve8 e850 (grid_evolve[850], grid[817], grid[818], grid[819], grid[849], grid[851], grid[881], grid[882], grid[883], grid[850]);
evolve8 e851 (grid_evolve[851], grid[818], grid[819], grid[820], grid[850], grid[852], grid[882], grid[883], grid[884], grid[851]);
evolve8 e852 (grid_evolve[852], grid[819], grid[820], grid[821], grid[851], grid[853], grid[883], grid[884], grid[885], grid[852]);
evolve8 e853 (grid_evolve[853], grid[820], grid[821], grid[822], grid[852], grid[854], grid[884], grid[885], grid[886], grid[853]);
evolve8 e854 (grid_evolve[854], grid[821], grid[822], grid[823], grid[853], grid[855], grid[885], grid[886], grid[887], grid[854]);
evolve8 e855 (grid_evolve[855], grid[822], grid[823], grid[824], grid[854], grid[856], grid[886], grid[887], grid[888], grid[855]);
evolve8 e856 (grid_evolve[856], grid[823], grid[824], grid[825], grid[855], grid[857], grid[887], grid[888], grid[889], grid[856]);
evolve8 e857 (grid_evolve[857], grid[824], grid[825], grid[826], grid[856], grid[858], grid[888], grid[889], grid[890], grid[857]);
evolve8 e858 (grid_evolve[858], grid[825], grid[826], grid[827], grid[857], grid[859], grid[889], grid[890], grid[891], grid[858]);
evolve8 e859 (grid_evolve[859], grid[826], grid[827], grid[828], grid[858], grid[860], grid[890], grid[891], grid[892], grid[859]);
evolve8 e860 (grid_evolve[860], grid[827], grid[828], grid[829], grid[859], grid[861], grid[891], grid[892], grid[893], grid[860]);
evolve8 e861 (grid_evolve[861], grid[828], grid[829], grid[830], grid[860], grid[862], grid[892], grid[893], grid[894], grid[861]);
evolve8 e862 (grid_evolve[862], grid[829], grid[830], grid[831], grid[861], grid[863], grid[893], grid[894], grid[895], grid[862]);
evolve5 e863 (grid_evolve[863], grid[830], grid[831], grid[862], grid[894], grid[895], grid[863]);

evolve5 e864 (grid_evolve[864], grid[832], grid[833], grid[865], grid[896], grid[897], grid[864]);
evolve8 e865 (grid_evolve[865], grid[832], grid[833], grid[834], grid[864], grid[866], grid[896], grid[897], grid[898], grid[865]);
evolve8 e866 (grid_evolve[866], grid[833], grid[834], grid[835], grid[865], grid[867], grid[897], grid[898], grid[899], grid[866]);
evolve8 e867 (grid_evolve[867], grid[834], grid[835], grid[836], grid[866], grid[868], grid[898], grid[899], grid[900], grid[867]);
evolve8 e868 (grid_evolve[868], grid[835], grid[836], grid[837], grid[867], grid[869], grid[899], grid[900], grid[901], grid[868]);
evolve8 e869 (grid_evolve[869], grid[836], grid[837], grid[838], grid[868], grid[870], grid[900], grid[901], grid[902], grid[869]);
evolve8 e870 (grid_evolve[870], grid[837], grid[838], grid[839], grid[869], grid[871], grid[901], grid[902], grid[903], grid[870]);
evolve8 e871 (grid_evolve[871], grid[838], grid[839], grid[840], grid[870], grid[872], grid[902], grid[903], grid[904], grid[871]);
evolve8 e872 (grid_evolve[872], grid[839], grid[840], grid[841], grid[871], grid[873], grid[903], grid[904], grid[905], grid[872]);
evolve8 e873 (grid_evolve[873], grid[840], grid[841], grid[842], grid[872], grid[874], grid[904], grid[905], grid[906], grid[873]);
evolve8 e874 (grid_evolve[874], grid[841], grid[842], grid[843], grid[873], grid[875], grid[905], grid[906], grid[907], grid[874]);
evolve8 e875 (grid_evolve[875], grid[842], grid[843], grid[844], grid[874], grid[876], grid[906], grid[907], grid[908], grid[875]);
evolve8 e876 (grid_evolve[876], grid[843], grid[844], grid[845], grid[875], grid[877], grid[907], grid[908], grid[909], grid[876]);
evolve8 e877 (grid_evolve[877], grid[844], grid[845], grid[846], grid[876], grid[878], grid[908], grid[909], grid[910], grid[877]);
evolve8 e878 (grid_evolve[878], grid[845], grid[846], grid[847], grid[877], grid[879], grid[909], grid[910], grid[911], grid[878]);
evolve8 e879 (grid_evolve[879], grid[846], grid[847], grid[848], grid[878], grid[880], grid[910], grid[911], grid[912], grid[879]);
evolve8 e880 (grid_evolve[880], grid[847], grid[848], grid[849], grid[879], grid[881], grid[911], grid[912], grid[913], grid[880]);
evolve8 e881 (grid_evolve[881], grid[848], grid[849], grid[850], grid[880], grid[882], grid[912], grid[913], grid[914], grid[881]);
evolve8 e882 (grid_evolve[882], grid[849], grid[850], grid[851], grid[881], grid[883], grid[913], grid[914], grid[915], grid[882]);
evolve8 e883 (grid_evolve[883], grid[850], grid[851], grid[852], grid[882], grid[884], grid[914], grid[915], grid[916], grid[883]);
evolve8 e884 (grid_evolve[884], grid[851], grid[852], grid[853], grid[883], grid[885], grid[915], grid[916], grid[917], grid[884]);
evolve8 e885 (grid_evolve[885], grid[852], grid[853], grid[854], grid[884], grid[886], grid[916], grid[917], grid[918], grid[885]);
evolve8 e886 (grid_evolve[886], grid[853], grid[854], grid[855], grid[885], grid[887], grid[917], grid[918], grid[919], grid[886]);
evolve8 e887 (grid_evolve[887], grid[854], grid[855], grid[856], grid[886], grid[888], grid[918], grid[919], grid[920], grid[887]);
evolve8 e888 (grid_evolve[888], grid[855], grid[856], grid[857], grid[887], grid[889], grid[919], grid[920], grid[921], grid[888]);
evolve8 e889 (grid_evolve[889], grid[856], grid[857], grid[858], grid[888], grid[890], grid[920], grid[921], grid[922], grid[889]);
evolve8 e890 (grid_evolve[890], grid[857], grid[858], grid[859], grid[889], grid[891], grid[921], grid[922], grid[923], grid[890]);
evolve8 e891 (grid_evolve[891], grid[858], grid[859], grid[860], grid[890], grid[892], grid[922], grid[923], grid[924], grid[891]);
evolve8 e892 (grid_evolve[892], grid[859], grid[860], grid[861], grid[891], grid[893], grid[923], grid[924], grid[925], grid[892]);
evolve8 e893 (grid_evolve[893], grid[860], grid[861], grid[862], grid[892], grid[894], grid[924], grid[925], grid[926], grid[893]);
evolve8 e894 (grid_evolve[894], grid[861], grid[862], grid[863], grid[893], grid[895], grid[925], grid[926], grid[927], grid[894]);
evolve5 e895 (grid_evolve[895], grid[862], grid[863], grid[894], grid[926], grid[927], grid[895]);

evolve5 e896 (grid_evolve[896], grid[864], grid[865], grid[897], grid[928], grid[929], grid[896]);
evolve8 e897 (grid_evolve[897], grid[864], grid[865], grid[866], grid[896], grid[898], grid[928], grid[929], grid[930], grid[897]);
evolve8 e898 (grid_evolve[898], grid[865], grid[866], grid[867], grid[897], grid[899], grid[929], grid[930], grid[931], grid[898]);
evolve8 e899 (grid_evolve[899], grid[866], grid[867], grid[868], grid[898], grid[900], grid[930], grid[931], grid[932], grid[899]);
evolve8 e900 (grid_evolve[900], grid[867], grid[868], grid[869], grid[899], grid[901], grid[931], grid[932], grid[933], grid[900]);
evolve8 e901 (grid_evolve[901], grid[868], grid[869], grid[870], grid[900], grid[902], grid[932], grid[933], grid[934], grid[901]);
evolve8 e902 (grid_evolve[902], grid[869], grid[870], grid[871], grid[901], grid[903], grid[933], grid[934], grid[935], grid[902]);
evolve8 e903 (grid_evolve[903], grid[870], grid[871], grid[872], grid[902], grid[904], grid[934], grid[935], grid[936], grid[903]);
evolve8 e904 (grid_evolve[904], grid[871], grid[872], grid[873], grid[903], grid[905], grid[935], grid[936], grid[937], grid[904]);
evolve8 e905 (grid_evolve[905], grid[872], grid[873], grid[874], grid[904], grid[906], grid[936], grid[937], grid[938], grid[905]);
evolve8 e906 (grid_evolve[906], grid[873], grid[874], grid[875], grid[905], grid[907], grid[937], grid[938], grid[939], grid[906]);
evolve8 e907 (grid_evolve[907], grid[874], grid[875], grid[876], grid[906], grid[908], grid[938], grid[939], grid[940], grid[907]);
evolve8 e908 (grid_evolve[908], grid[875], grid[876], grid[877], grid[907], grid[909], grid[939], grid[940], grid[941], grid[908]);
evolve8 e909 (grid_evolve[909], grid[876], grid[877], grid[878], grid[908], grid[910], grid[940], grid[941], grid[942], grid[909]);
evolve8 e910 (grid_evolve[910], grid[877], grid[878], grid[879], grid[909], grid[911], grid[941], grid[942], grid[943], grid[910]);
evolve8 e911 (grid_evolve[911], grid[878], grid[879], grid[880], grid[910], grid[912], grid[942], grid[943], grid[944], grid[911]);
evolve8 e912 (grid_evolve[912], grid[879], grid[880], grid[881], grid[911], grid[913], grid[943], grid[944], grid[945], grid[912]);
evolve8 e913 (grid_evolve[913], grid[880], grid[881], grid[882], grid[912], grid[914], grid[944], grid[945], grid[946], grid[913]);
evolve8 e914 (grid_evolve[914], grid[881], grid[882], grid[883], grid[913], grid[915], grid[945], grid[946], grid[947], grid[914]);
evolve8 e915 (grid_evolve[915], grid[882], grid[883], grid[884], grid[914], grid[916], grid[946], grid[947], grid[948], grid[915]);
evolve8 e916 (grid_evolve[916], grid[883], grid[884], grid[885], grid[915], grid[917], grid[947], grid[948], grid[949], grid[916]);
evolve8 e917 (grid_evolve[917], grid[884], grid[885], grid[886], grid[916], grid[918], grid[948], grid[949], grid[950], grid[917]);
evolve8 e918 (grid_evolve[918], grid[885], grid[886], grid[887], grid[917], grid[919], grid[949], grid[950], grid[951], grid[918]);
evolve8 e919 (grid_evolve[919], grid[886], grid[887], grid[888], grid[918], grid[920], grid[950], grid[951], grid[952], grid[919]);
evolve8 e920 (grid_evolve[920], grid[887], grid[888], grid[889], grid[919], grid[921], grid[951], grid[952], grid[953], grid[920]);
evolve8 e921 (grid_evolve[921], grid[888], grid[889], grid[890], grid[920], grid[922], grid[952], grid[953], grid[954], grid[921]);
evolve8 e922 (grid_evolve[922], grid[889], grid[890], grid[891], grid[921], grid[923], grid[953], grid[954], grid[955], grid[922]);
evolve8 e923 (grid_evolve[923], grid[890], grid[891], grid[892], grid[922], grid[924], grid[954], grid[955], grid[956], grid[923]);
evolve8 e924 (grid_evolve[924], grid[891], grid[892], grid[893], grid[923], grid[925], grid[955], grid[956], grid[957], grid[924]);
evolve8 e925 (grid_evolve[925], grid[892], grid[893], grid[894], grid[924], grid[926], grid[956], grid[957], grid[958], grid[925]);
evolve8 e926 (grid_evolve[926], grid[893], grid[894], grid[895], grid[925], grid[927], grid[957], grid[958], grid[959], grid[926]);
evolve5 e927 (grid_evolve[927], grid[894], grid[895], grid[926], grid[958], grid[959], grid[927]);

evolve5 e928 (grid_evolve[928], grid[896], grid[897], grid[929], grid[960], grid[961], grid[928]);
evolve8 e929 (grid_evolve[929], grid[896], grid[897], grid[898], grid[928], grid[930], grid[960], grid[961], grid[962], grid[929]);
evolve8 e930 (grid_evolve[930], grid[897], grid[898], grid[899], grid[929], grid[931], grid[961], grid[962], grid[963], grid[930]);
evolve8 e931 (grid_evolve[931], grid[898], grid[899], grid[900], grid[930], grid[932], grid[962], grid[963], grid[964], grid[931]);
evolve8 e932 (grid_evolve[932], grid[899], grid[900], grid[901], grid[931], grid[933], grid[963], grid[964], grid[965], grid[932]);
evolve8 e933 (grid_evolve[933], grid[900], grid[901], grid[902], grid[932], grid[934], grid[964], grid[965], grid[966], grid[933]);
evolve8 e934 (grid_evolve[934], grid[901], grid[902], grid[903], grid[933], grid[935], grid[965], grid[966], grid[967], grid[934]);
evolve8 e935 (grid_evolve[935], grid[902], grid[903], grid[904], grid[934], grid[936], grid[966], grid[967], grid[968], grid[935]);
evolve8 e936 (grid_evolve[936], grid[903], grid[904], grid[905], grid[935], grid[937], grid[967], grid[968], grid[969], grid[936]);
evolve8 e937 (grid_evolve[937], grid[904], grid[905], grid[906], grid[936], grid[938], grid[968], grid[969], grid[970], grid[937]);
evolve8 e938 (grid_evolve[938], grid[905], grid[906], grid[907], grid[937], grid[939], grid[969], grid[970], grid[971], grid[938]);
evolve8 e939 (grid_evolve[939], grid[906], grid[907], grid[908], grid[938], grid[940], grid[970], grid[971], grid[972], grid[939]);
evolve8 e940 (grid_evolve[940], grid[907], grid[908], grid[909], grid[939], grid[941], grid[971], grid[972], grid[973], grid[940]);
evolve8 e941 (grid_evolve[941], grid[908], grid[909], grid[910], grid[940], grid[942], grid[972], grid[973], grid[974], grid[941]);
evolve8 e942 (grid_evolve[942], grid[909], grid[910], grid[911], grid[941], grid[943], grid[973], grid[974], grid[975], grid[942]);
evolve8 e943 (grid_evolve[943], grid[910], grid[911], grid[912], grid[942], grid[944], grid[974], grid[975], grid[976], grid[943]);
evolve8 e944 (grid_evolve[944], grid[911], grid[912], grid[913], grid[943], grid[945], grid[975], grid[976], grid[977], grid[944]);
evolve8 e945 (grid_evolve[945], grid[912], grid[913], grid[914], grid[944], grid[946], grid[976], grid[977], grid[978], grid[945]);
evolve8 e946 (grid_evolve[946], grid[913], grid[914], grid[915], grid[945], grid[947], grid[977], grid[978], grid[979], grid[946]);
evolve8 e947 (grid_evolve[947], grid[914], grid[915], grid[916], grid[946], grid[948], grid[978], grid[979], grid[980], grid[947]);
evolve8 e948 (grid_evolve[948], grid[915], grid[916], grid[917], grid[947], grid[949], grid[979], grid[980], grid[981], grid[948]);
evolve8 e949 (grid_evolve[949], grid[916], grid[917], grid[918], grid[948], grid[950], grid[980], grid[981], grid[982], grid[949]);
evolve8 e950 (grid_evolve[950], grid[917], grid[918], grid[919], grid[949], grid[951], grid[981], grid[982], grid[983], grid[950]);
evolve8 e951 (grid_evolve[951], grid[918], grid[919], grid[920], grid[950], grid[952], grid[982], grid[983], grid[984], grid[951]);
evolve8 e952 (grid_evolve[952], grid[919], grid[920], grid[921], grid[951], grid[953], grid[983], grid[984], grid[985], grid[952]);
evolve8 e953 (grid_evolve[953], grid[920], grid[921], grid[922], grid[952], grid[954], grid[984], grid[985], grid[986], grid[953]);
evolve8 e954 (grid_evolve[954], grid[921], grid[922], grid[923], grid[953], grid[955], grid[985], grid[986], grid[987], grid[954]);
evolve8 e955 (grid_evolve[955], grid[922], grid[923], grid[924], grid[954], grid[956], grid[986], grid[987], grid[988], grid[955]);
evolve8 e956 (grid_evolve[956], grid[923], grid[924], grid[925], grid[955], grid[957], grid[987], grid[988], grid[989], grid[956]);
evolve8 e957 (grid_evolve[957], grid[924], grid[925], grid[926], grid[956], grid[958], grid[988], grid[989], grid[990], grid[957]);
evolve8 e958 (grid_evolve[958], grid[925], grid[926], grid[927], grid[957], grid[959], grid[989], grid[990], grid[991], grid[958]);
evolve5 e959 (grid_evolve[959], grid[926], grid[927], grid[958], grid[990], grid[991], grid[959]);

evolve5 e960 (grid_evolve[960], grid[928], grid[929], grid[961], grid[992], grid[993], grid[960]);
evolve8 e961 (grid_evolve[961], grid[928], grid[929], grid[930], grid[960], grid[962], grid[992], grid[993], grid[994], grid[961]);
evolve8 e962 (grid_evolve[962], grid[929], grid[930], grid[931], grid[961], grid[963], grid[993], grid[994], grid[995], grid[962]);
evolve8 e963 (grid_evolve[963], grid[930], grid[931], grid[932], grid[962], grid[964], grid[994], grid[995], grid[996], grid[963]);
evolve8 e964 (grid_evolve[964], grid[931], grid[932], grid[933], grid[963], grid[965], grid[995], grid[996], grid[997], grid[964]);
evolve8 e965 (grid_evolve[965], grid[932], grid[933], grid[934], grid[964], grid[966], grid[996], grid[997], grid[998], grid[965]);
evolve8 e966 (grid_evolve[966], grid[933], grid[934], grid[935], grid[965], grid[967], grid[997], grid[998], grid[999], grid[966]);
evolve8 e967 (grid_evolve[967], grid[934], grid[935], grid[936], grid[966], grid[968], grid[998], grid[999], grid[1000], grid[967]);
evolve8 e968 (grid_evolve[968], grid[935], grid[936], grid[937], grid[967], grid[969], grid[999], grid[1000], grid[1001], grid[968]);
evolve8 e969 (grid_evolve[969], grid[936], grid[937], grid[938], grid[968], grid[970], grid[1000], grid[1001], grid[1002], grid[969]);
evolve8 e970 (grid_evolve[970], grid[937], grid[938], grid[939], grid[969], grid[971], grid[1001], grid[1002], grid[1003], grid[970]);
evolve8 e971 (grid_evolve[971], grid[938], grid[939], grid[940], grid[970], grid[972], grid[1002], grid[1003], grid[1004], grid[971]);
evolve8 e972 (grid_evolve[972], grid[939], grid[940], grid[941], grid[971], grid[973], grid[1003], grid[1004], grid[1005], grid[972]);
evolve8 e973 (grid_evolve[973], grid[940], grid[941], grid[942], grid[972], grid[974], grid[1004], grid[1005], grid[1006], grid[973]);
evolve8 e974 (grid_evolve[974], grid[941], grid[942], grid[943], grid[973], grid[975], grid[1005], grid[1006], grid[1007], grid[974]);
evolve8 e975 (grid_evolve[975], grid[942], grid[943], grid[944], grid[974], grid[976], grid[1006], grid[1007], grid[1008], grid[975]);
evolve8 e976 (grid_evolve[976], grid[943], grid[944], grid[945], grid[975], grid[977], grid[1007], grid[1008], grid[1009], grid[976]);
evolve8 e977 (grid_evolve[977], grid[944], grid[945], grid[946], grid[976], grid[978], grid[1008], grid[1009], grid[1010], grid[977]);
evolve8 e978 (grid_evolve[978], grid[945], grid[946], grid[947], grid[977], grid[979], grid[1009], grid[1010], grid[1011], grid[978]);
evolve8 e979 (grid_evolve[979], grid[946], grid[947], grid[948], grid[978], grid[980], grid[1010], grid[1011], grid[1012], grid[979]);
evolve8 e980 (grid_evolve[980], grid[947], grid[948], grid[949], grid[979], grid[981], grid[1011], grid[1012], grid[1013], grid[980]);
evolve8 e981 (grid_evolve[981], grid[948], grid[949], grid[950], grid[980], grid[982], grid[1012], grid[1013], grid[1014], grid[981]);
evolve8 e982 (grid_evolve[982], grid[949], grid[950], grid[951], grid[981], grid[983], grid[1013], grid[1014], grid[1015], grid[982]);
evolve8 e983 (grid_evolve[983], grid[950], grid[951], grid[952], grid[982], grid[984], grid[1014], grid[1015], grid[1016], grid[983]);
evolve8 e984 (grid_evolve[984], grid[951], grid[952], grid[953], grid[983], grid[985], grid[1015], grid[1016], grid[1017], grid[984]);
evolve8 e985 (grid_evolve[985], grid[952], grid[953], grid[954], grid[984], grid[986], grid[1016], grid[1017], grid[1018], grid[985]);
evolve8 e986 (grid_evolve[986], grid[953], grid[954], grid[955], grid[985], grid[987], grid[1017], grid[1018], grid[1019], grid[986]);
evolve8 e987 (grid_evolve[987], grid[954], grid[955], grid[956], grid[986], grid[988], grid[1018], grid[1019], grid[1020], grid[987]);
evolve8 e988 (grid_evolve[988], grid[955], grid[956], grid[957], grid[987], grid[989], grid[1019], grid[1020], grid[1021], grid[988]);
evolve8 e989 (grid_evolve[989], grid[956], grid[957], grid[958], grid[988], grid[990], grid[1020], grid[1021], grid[1022], grid[989]);
evolve8 e990 (grid_evolve[990], grid[957], grid[958], grid[959], grid[989], grid[991], grid[1021], grid[1022], grid[1023], grid[990]);
evolve5 e991 (grid_evolve[991], grid[958], grid[959], grid[990], grid[1022], grid[1023], grid[991]);

evolve3 e992 (grid_evolve[992], grid[960], grid[961], grid[993], grid[992]);
evolve5 e993 (grid_evolve[993], grid[960], grid[961], grid[962], grid[992], grid[994], grid[993]);
evolve5 e994 (grid_evolve[994], grid[961], grid[962], grid[963], grid[993], grid[995], grid[994]);
evolve5 e995 (grid_evolve[995], grid[962], grid[963], grid[964], grid[994], grid[996], grid[995]);
evolve5 e996 (grid_evolve[996], grid[963], grid[964], grid[965], grid[995], grid[997], grid[996]);
evolve5 e997 (grid_evolve[997], grid[964], grid[965], grid[966], grid[996], grid[998], grid[997]);
evolve5 e998 (grid_evolve[998], grid[965], grid[966], grid[967], grid[997], grid[999], grid[998]);
evolve5 e999 (grid_evolve[999], grid[966], grid[967], grid[968], grid[998], grid[1000], grid[999]);
evolve5 e1000 (grid_evolve[1000], grid[967], grid[968], grid[969], grid[999], grid[1001], grid[1000]);
evolve5 e1001 (grid_evolve[1001], grid[968], grid[969], grid[970], grid[1000], grid[1002], grid[1001]);
evolve5 e1002 (grid_evolve[1002], grid[969], grid[970], grid[971], grid[1001], grid[1003], grid[1002]);
evolve5 e1003 (grid_evolve[1003], grid[970], grid[971], grid[972], grid[1002], grid[1004], grid[1003]);
evolve5 e1004 (grid_evolve[1004], grid[971], grid[972], grid[973], grid[1003], grid[1005], grid[1004]);
evolve5 e1005 (grid_evolve[1005], grid[972], grid[973], grid[974], grid[1004], grid[1006], grid[1005]);
evolve5 e1006 (grid_evolve[1006], grid[973], grid[974], grid[975], grid[1005], grid[1007], grid[1006]);
evolve5 e1007 (grid_evolve[1007], grid[974], grid[975], grid[976], grid[1006], grid[1008], grid[1007]);
evolve5 e1008 (grid_evolve[1008], grid[975], grid[976], grid[977], grid[1007], grid[1009], grid[1008]);
evolve5 e1009 (grid_evolve[1009], grid[976], grid[977], grid[978], grid[1008], grid[1010], grid[1009]);
evolve5 e1010 (grid_evolve[1010], grid[977], grid[978], grid[979], grid[1009], grid[1011], grid[1010]);
evolve5 e1011 (grid_evolve[1011], grid[978], grid[979], grid[980], grid[1010], grid[1012], grid[1011]);
evolve5 e1012 (grid_evolve[1012], grid[979], grid[980], grid[981], grid[1011], grid[1013], grid[1012]);
evolve5 e1013 (grid_evolve[1013], grid[980], grid[981], grid[982], grid[1012], grid[1014], grid[1013]);
evolve5 e1014 (grid_evolve[1014], grid[981], grid[982], grid[983], grid[1013], grid[1015], grid[1014]);
evolve5 e1015 (grid_evolve[1015], grid[982], grid[983], grid[984], grid[1014], grid[1016], grid[1015]);
evolve5 e1016 (grid_evolve[1016], grid[983], grid[984], grid[985], grid[1015], grid[1017], grid[1016]);
evolve5 e1017 (grid_evolve[1017], grid[984], grid[985], grid[986], grid[1016], grid[1018], grid[1017]);
evolve5 e1018 (grid_evolve[1018], grid[985], grid[986], grid[987], grid[1017], grid[1019], grid[1018]);
evolve5 e1019 (grid_evolve[1019], grid[986], grid[987], grid[988], grid[1018], grid[1020], grid[1019]);
evolve5 e1020 (grid_evolve[1020], grid[987], grid[988], grid[989], grid[1019], grid[1021], grid[1020]);
evolve5 e1021 (grid_evolve[1021], grid[988], grid[989], grid[990], grid[1020], grid[1022], grid[1021]);
evolve5 e1022 (grid_evolve[1022], grid[989], grid[990], grid[991], grid[1021], grid[1023], grid[1022]);
evolve3 e1023 (grid_evolve[1023], grid[990], grid[991], grid[1022], grid[1023]);



endmodule // top


module evolve3 (next_state, vector1, vector2, vector3, current_state);
	
   input logic  vector1;
   input logic  vector2;
   input logic  vector3;
   input logic  current_state;
   output logic next_state;
   
   logic [3:0] 	sum;
   
   assign sum = vector1 + vector2 + vector3;
   rules r1 (sum, current_state, next_state);
   
endmodule // evolve3

module evolve5 (next_state, vector1, vector2, vector3, 
		vector4, vector5, current_state);
   
   input logic   vector1;
   input logic 	 vector2;
   input logic 	 vector3;
   input logic 	 vector4;
   input logic 	 vector5;
   input logic 	 current_state;
   output logic  next_state;
   
   logic [3:0] 	 sum;
   
   assign sum = vector1 + vector2 + vector3 + vector4 + vector5;
   rules r1 (sum, current_state, next_state);
   
endmodule // evolve5


module evolve8 (next_state, vector1, vector2, vector3, 
		vector4, vector5, vector6, 
		vector7, vector8, current_state);
   
   input logic 	vector1;
   input logic 	vector2;
   input logic 	vector3;
   input logic 	vector4;
   input logic 	vector5;
	
   input logic 	vector6;
   input logic 	vector7;
   input logic 	vector8;
   input logic 	current_state;
   output logic next_state;
   
   logic [3:0] 	sum;
   
   assign sum = vector1 + vector2 + vector3 + vector4 + 
		vector5 + vector6 + vector7 + vector8;
   rules r1 (sum, current_state, next_state);
   
endmodule // evolve8


module rules (pop_count, current_state, next_state);
   
   input logic [3:0] pop_count;
   input logic 	     current_state;
   output logic      next_state;
   
   assign next_state = (pop_count == 2 & current_state) | pop_count == 3;
   
endmodule // rules





